`timescale 1ns/1ps

module tb_polymult();
    // Parameters
    parameter WORD_WIDTH = 32;
    parameter MEM_SIZE = 553;
    parameter MEM_SPARSE_SIZE = 50;
    parameter CLK_PERIOD = 10;

    // Test data - Normal words array
    reg [WORD_WIDTH-1:0] normal_words [0:MEM_SIZE - 1];
    reg [WORD_WIDTH-1:0] acc_words [0:MEM_SIZE - 1];
    
    // Sparse memory data pairs
    reg [31:0] sparse_pairs [0:MEM_SPARSE_SIZE-1];

    // Signals
    reg clk;
    reg rst_n;
    reg [WORD_WIDTH-1:0] normal_mem_data_i;
    reg [WORD_WIDTH-1:0] sparse_mem_data_i;
    reg [WORD_WIDTH-1:0] acc_mem_data_i;
    reg [9:0] sparse_mem_addr_i;
    reg start_process;

    reg [9:0] acc_start_idx_high;
    reg [9:0] acc_start_idx_low;
    reg [4:0] high_low_diff;


    wire [WORD_WIDTH-1:0] acc_mem_write_data_o;
    wire acc_mem_write_en;
    wire [9:0] normal_mem_addr_o;
    wire [9:0] acc_mem_addr_o;
    wire process_done;
    wire busy;

    // Clock generation
    initial begin
        clk = 0;
        forever #(CLK_PERIOD/2) clk = ~clk;
    end

    // Declare integer for loop iteration
    integer i;
    integer pair_idx;
    integer word_index;
    integer bit_index;


    // Declare bit_positions array
    


    // DUT instantiation
    controller #(
        .WORD_WIDTH(WORD_WIDTH),
        .MEM_SIZE(MEM_SIZE),
        .MEM_SPARSE_SIZE(MEM_SPARSE_SIZE)
    ) dut (
        .clk(clk),
        .rst_n(rst_n),
        .normal_mem_data_i(normal_mem_data_i),
        .sparse_mem_data_i(sparse_mem_data_i),
        .acc_mem_data_i(acc_mem_data_i),
        .sparse_mem_addr_i(sparse_mem_addr_i),
        .acc_mem_write_data_o(acc_mem_write_data_o),
        .acc_mem_write_en(acc_mem_write_en),
        .normal_mem_addr_o(normal_mem_addr_o),
        .acc_mem_addr_o(acc_mem_addr_o),
        .start_process(start_process),
        .process_done(process_done),
        .busy(busy)
    );

    // Test stimulus
    initial begin
        // Initialize inputs
        for(i = 0; i < MEM_SIZE; i = i + 1) begin
            acc_words[i] = 32'b0;
            normal_words[i] = 32'b0;
        end


        normal_words[0] = 32'b11110110000000010101100010011100;
        normal_words[1] = 32'b00110011111110101100111000011011;
        normal_words[2] = 32'b00100011001100100011100011101001;
        normal_words[3] = 32'b00011010000010100001000101100000;
        normal_words[4] = 32'b11111101011111011010010100110110;
        normal_words[5] = 32'b10001101011010101100111010101101;
        normal_words[6] = 32'b10111111100000000101011110000111;
        normal_words[7] = 32'b11001001100110011011011100100101;
        normal_words[8] = 32'b01000000110100010011110111011011;
        normal_words[9] = 32'b00100101101110010000010101100110;
        normal_words[10] = 32'b00100111100111111100110001001100;
        normal_words[11] = 32'b10111010100110010001101000111101;
        normal_words[12] = 32'b10010000111100111001000001111001;
        normal_words[13] = 32'b01001110011110100110110001101101;
        normal_words[14] = 32'b11101011000000110011101100010000;
        normal_words[15] = 32'b01100110101010000101100111111101;
        normal_words[16] = 32'b00011110101100110011001000110110;
        normal_words[17] = 32'b01011101100000011010110010101010;
        normal_words[18] = 32'b01000000001110011011111010000100;
        normal_words[19] = 32'b01011011010110101000001100010110;
        normal_words[20] = 32'b00110100000101100010110101011001;
        normal_words[21] = 32'b11011000011110001110011101001110;
        normal_words[22] = 32'b01011101001011011010101101001001;
        normal_words[23] = 32'b10110100011011111000011000111111;
        normal_words[24] = 32'b00101101001100010000101110001011;
        normal_words[25] = 32'b01111001001011100010001000000110;
        normal_words[26] = 32'b01111010101110101001100011100101;
        normal_words[27] = 32'b01111001111011111001110010101001;
        normal_words[28] = 32'b11011101011100000001001111100000;
        normal_words[29] = 32'b00111111101110000000100111111011;
        normal_words[30] = 32'b10111101010110100000110011101101;
        normal_words[31] = 32'b00101011000010011011111111000000;
        normal_words[32] = 32'b11011101011001001100111010011100;
        normal_words[33] = 32'b11111001100011101000000001110010;
        normal_words[34] = 32'b01011110111011011000101001010000;
        normal_words[35] = 32'b10010111011000010110010101001001;
        normal_words[36] = 32'b00001010101000010010001101111011;
        normal_words[37] = 32'b00111101100101111100110110110010;
        normal_words[38] = 32'b10011000011110011111110011010101;
        normal_words[39] = 32'b11100110010111110001010111001010;
        normal_words[40] = 32'b10011111101111101110011001111101;
        normal_words[41] = 32'b01111011110011110100001010010110;
        normal_words[42] = 32'b11010000100010101111010011001110;
        normal_words[43] = 32'b10011110001000011011001010101011;
        normal_words[44] = 32'b10110110111100001000011110010001;
        normal_words[45] = 32'b10110000101001101011001110000111;
        normal_words[46] = 32'b01101100001111011111111101001000;
        normal_words[47] = 32'b11100000100111001111011011111110;
        normal_words[48] = 32'b10111000010010100111101101000100;
        normal_words[49] = 32'b00110100101100000110000111011011;
        normal_words[50] = 32'b10100101001010101011010100111101;
        normal_words[51] = 32'b00101110111000000101111111000111;
        normal_words[52] = 32'b10101101100011011111010100110110;
        normal_words[53] = 32'b11100001110000011110000110101110;
        normal_words[54] = 32'b11011000011000010010000000000001;
        normal_words[55] = 32'b10100010100011011000111100001110;
        normal_words[56] = 32'b00010101101011100111001010110011;
        normal_words[57] = 32'b10010100101001010111001111100010;
        normal_words[58] = 32'b00101110011000111100101011011011;
        normal_words[59] = 32'b01101101001111101010100111000011;
        normal_words[60] = 32'b00000001000101010011110001010111;
        normal_words[61] = 32'b11101100000110011001011101011110;
        normal_words[62] = 32'b10011101010110010000101101111010;
        normal_words[63] = 32'b01001010001110100101111110110101;
        normal_words[64] = 32'b01011001011011111111000001111110;
        normal_words[65] = 32'b10100011101011100101010111110110;
        normal_words[66] = 32'b01000100101000101011110110111111;
        normal_words[67] = 32'b11110011110011110111111101001011;
        normal_words[68] = 32'b11100100011111110001000010100111;
        normal_words[69] = 32'b11011100001000100000100100110101;
        normal_words[70] = 32'b00101101001111110110010101001100;
        normal_words[71] = 32'b00000111001011101011110110110100;
        normal_words[72] = 32'b11011010001011001010010100100111;
        normal_words[73] = 32'b10000101000011101010101111100001;
        normal_words[74] = 32'b00110100101100101111110100011110;
        normal_words[75] = 32'b11101101101001000110000111111110;
        normal_words[76] = 32'b01101111011000001100101001110101;
        normal_words[77] = 32'b01001100000111111011100001110101;
        normal_words[78] = 32'b11101010010011101000101110010011;
        normal_words[79] = 32'b00111001000000001010100111000110;
        normal_words[80] = 32'b00111101100111111011000101111000;
        normal_words[81] = 32'b11010110111110100011101000111111;
        normal_words[82] = 32'b01100000000110001001111100001011;
        normal_words[83] = 32'b10000001010011010001110100000111;
        normal_words[84] = 32'b10010101110010000110001111100110;
        normal_words[85] = 32'b00100101100110101110000100111000;
        normal_words[86] = 32'b11010101011011101000110111110000;
        normal_words[87] = 32'b11110110010100000001000001011111;
        normal_words[88] = 32'b00010011100100101101011000111111;
        normal_words[89] = 32'b00000111010101000100000111100101;
        normal_words[90] = 32'b00010100011010111010110011000101;
        normal_words[91] = 32'b10001001000001111011111100010100;
        normal_words[92] = 32'b10100111110000110100011111110000;
        normal_words[93] = 32'b10011010110000001111111101100011;
        normal_words[94] = 32'b11100001001101010100000100001010;
        normal_words[95] = 32'b11001011111110110100001001010001;
        normal_words[96] = 32'b10101010001000100010000101101100;
        normal_words[97] = 32'b11001011111110001100010101010101;
        normal_words[98] = 32'b11100011111000011001110111011100;
        normal_words[99] = 32'b10010100011011001100101101101101;
        normal_words[100] = 32'b00111011100101101111000011001101;
        normal_words[101] = 32'b00000110101101110110100101101110;
        normal_words[102] = 32'b01101110101101101111111100010000;
        normal_words[103] = 32'b01110000111101000101101111010011;
        normal_words[104] = 32'b11101101011100101101111001100101;
        normal_words[105] = 32'b00100100001010111100000100111010;
        normal_words[106] = 32'b10101001001101110000110110001000;
        normal_words[107] = 32'b01001010000111100110000000010110;
        normal_words[108] = 32'b11011011110010010110110000000011;
        normal_words[109] = 32'b11101011011111110000000000101011;
        normal_words[110] = 32'b11100110110001000111010011111100;
        normal_words[111] = 32'b11000100010100000001111011100101;
        normal_words[112] = 32'b11010011011111010100101010000111;
        normal_words[113] = 32'b10110000010101100001001001011011;
        normal_words[114] = 32'b00111100100011011010101001000100;
        normal_words[115] = 32'b00111001010101001001010110000000;
        normal_words[116] = 32'b10001001001110000111011010111111;
        normal_words[117] = 32'b11000111001011101101001101101011;
        normal_words[118] = 32'b00011100101111101000110100010110;
        normal_words[119] = 32'b10110000100010100111111101101111;
        normal_words[120] = 32'b11010100001000001100110011010010;
        normal_words[121] = 32'b00001010000011001010000111010110;
        normal_words[122] = 32'b01111011111101101110011011100111;
        normal_words[123] = 32'b11110110101100011110000000001011;
        normal_words[124] = 32'b01001111001101010010101000000110;
        normal_words[125] = 32'b00000101011100011110110001010101;
        normal_words[126] = 32'b10110111001001000111101001111111;
        normal_words[127] = 32'b10100010011110111010110101011001;
        normal_words[128] = 32'b00010010100001000001000010101111;
        normal_words[129] = 32'b11011111010010011000100011110111;
        normal_words[130] = 32'b10101100110111111101001010111111;
        normal_words[131] = 32'b10110010001111000000010110110101;
        normal_words[132] = 32'b10011111001100010001000010110011;
        normal_words[133] = 32'b11011010111011101010011000001100;
        normal_words[134] = 32'b01111000001000101010110010100001;
        normal_words[135] = 32'b10110100100111010100010110100011;
        normal_words[136] = 32'b11011001011111010000011101101100;
        normal_words[137] = 32'b00010100110110000110001100001110;
        normal_words[138] = 32'b11110100000010011110001101011010;
        normal_words[139] = 32'b00111000001101000010011001011010;
        normal_words[140] = 32'b11000011110010100111011000110010;
        normal_words[141] = 32'b00110000110110100000010011010101;
        normal_words[142] = 32'b00100010110010100010001011001001;
        normal_words[143] = 32'b10101101011000111100101010010111;
        normal_words[144] = 32'b00101001101111001011011111110011;
        normal_words[145] = 32'b10001111100000101100001100111100;
        normal_words[146] = 32'b10110000100111101001101100100101;
        normal_words[147] = 32'b01010101111111011110110111101011;
        normal_words[148] = 32'b01011010000001100100111011000000;
        normal_words[149] = 32'b10000000101101000001010110010100;
        normal_words[150] = 32'b11001000100001001111011000100100;
        normal_words[151] = 32'b01010100011000001100111001010010;
        normal_words[152] = 32'b10010110010111011111111010001111;
        normal_words[153] = 32'b10011001000101011010010011100001;
        normal_words[154] = 32'b01111001101101111111111000101100;
        normal_words[155] = 32'b01100111010011110011111001110101;
        normal_words[156] = 32'b10100101101010110100001001000001;
        normal_words[157] = 32'b10000111111010000101110111010110;
        normal_words[158] = 32'b00011001100000011000101111000000;
        normal_words[159] = 32'b00111010001010111100110010101011;
        normal_words[160] = 32'b10100111001010010000000101000100;
        normal_words[161] = 32'b01111101111010010011001001110011;
        normal_words[162] = 32'b01100101111001110100111110110100;
        normal_words[163] = 32'b10001100110000101100011000011011;
        normal_words[164] = 32'b00101101111011110011001000010011;
        normal_words[165] = 32'b10001110000101100111011010011111;
        normal_words[166] = 32'b11111100100001110101111001111110;
        normal_words[167] = 32'b11100111111110011101001001001111;
        normal_words[168] = 32'b10110001011101010110000001111101;
        normal_words[169] = 32'b00111011100111010010110001110101;
        normal_words[170] = 32'b10011110010101011111111111011110;
        normal_words[171] = 32'b11001101110010011011100010110110;
        normal_words[172] = 32'b01111110101010000001111100000001;
        normal_words[173] = 32'b11101000011001111000000101010100;
        normal_words[174] = 32'b11110101110101101011111011100000;
        normal_words[175] = 32'b01101100011111001001001011110101;
        normal_words[176] = 32'b10101010001100010010100011111111;
        normal_words[177] = 32'b01110010110100111011100110000001;
        normal_words[178] = 32'b00100001100101100100010001110110;
        normal_words[179] = 32'b00101101001101010101110010100110;
        normal_words[180] = 32'b10010000101110010001110011100000;
        normal_words[181] = 32'b00010101001010011010001100100000;
        normal_words[182] = 32'b11001011100000101100111010100001;
        normal_words[183] = 32'b01001101111001010100011100000100;
        normal_words[184] = 32'b00010000101111110000110101001111;
        normal_words[185] = 32'b01011101011101111110011011001011;
        normal_words[186] = 32'b10011111011010001001111001101011;
        normal_words[187] = 32'b11110010101111000011001011010011;
        normal_words[188] = 32'b11110011000100110100100100011101;
        normal_words[189] = 32'b11010100000100001001101011101111;
        normal_words[190] = 32'b11000100011001011100110111110011;
        normal_words[191] = 32'b00001110010001010001101001110111;
        normal_words[192] = 32'b10110110011111011110110111110101;
        normal_words[193] = 32'b01000101101111010101000101100011;
        normal_words[194] = 32'b01011011100010001101110111110110;
        normal_words[195] = 32'b00101100000101001110110100100100;
        normal_words[196] = 32'b01010011100110001101000110111011;
        normal_words[197] = 32'b01000010110101011010000000011100;
        normal_words[198] = 32'b11110000011001000110100101000110;
        normal_words[199] = 32'b01101100111000110111010111111001;
        normal_words[200] = 32'b00000010000111110010101001000110;
        normal_words[201] = 32'b00110111101010010111000110100100;
        normal_words[202] = 32'b10000010100111100101010011100011;
        normal_words[203] = 32'b11001000010001010000101011000110;
        normal_words[204] = 32'b10101011101000111110010001101010;
        normal_words[205] = 32'b10101010111000011100000011111111;
        normal_words[206] = 32'b10100101001011111010000011100010;
        normal_words[207] = 32'b00001001110001011010011111011111;
        normal_words[208] = 32'b00001110101000001110000010101110;
        normal_words[209] = 32'b11100111111100011111000011001111;
        normal_words[210] = 32'b11010010100000110000101100111000;
        normal_words[211] = 32'b11010001010110100001000101111010;
        normal_words[212] = 32'b01101100111010011000011000010001;
        normal_words[213] = 32'b11000001011111010000001011011010;
        normal_words[214] = 32'b10010011011011000111011001011110;
        normal_words[215] = 32'b00100010110000100000110100101001;
        normal_words[216] = 32'b01111001000000001010010000101100;
        normal_words[217] = 32'b01011110010011011001010001101111;
        normal_words[218] = 32'b10111100110001001110101101101001;
        normal_words[219] = 32'b00100000111001001111101001101101;
        normal_words[220] = 32'b01001001010110100111100001011100;
        normal_words[221] = 32'b10111110011001010101001010111111;
        normal_words[222] = 32'b01100110100000101101101011010000;
        normal_words[223] = 32'b00110011100101011010100101101110;
        normal_words[224] = 32'b10001110110110111101110100101110;
        normal_words[225] = 32'b01100110101011100010100100011001;
        normal_words[226] = 32'b00010001001000010101100001001010;
        normal_words[227] = 32'b11111010111000000010111010111110;
        normal_words[228] = 32'b11100110011100010110111011111011;
        normal_words[229] = 32'b10011010100000000011011110101110;
        normal_words[230] = 32'b01100001011000110010000111111001;
        normal_words[231] = 32'b01010010000000010011001000111000;
        normal_words[232] = 32'b00000111000111100011011000010011;
        normal_words[233] = 32'b11001011001101101000011110001010;
        normal_words[234] = 32'b00110001001000110101111110100110;
        normal_words[235] = 32'b10001011110111010000101101001000;
        normal_words[236] = 32'b01101101001111111111111001100001;
        normal_words[237] = 32'b11111000110111001011111101101000;
        normal_words[238] = 32'b00000011101001001000001001101110;
        normal_words[239] = 32'b10011100100010110101101010100101;
        normal_words[240] = 32'b10100011011001011011000001001111;
        normal_words[241] = 32'b11101111101110110100001101100010;
        normal_words[242] = 32'b00101111101011110001011000100000;
        normal_words[243] = 32'b10100101101111100010000111111111;
        normal_words[244] = 32'b00010101001101011001010101011010;
        normal_words[245] = 32'b01110111110000101011111000001000;
        normal_words[246] = 32'b01010110001111001011100101101011;
        normal_words[247] = 32'b10111001001000001101101000100101;
        normal_words[248] = 32'b01111100110001011110110000101111;
        normal_words[249] = 32'b00001000001000001110001010001011;
        normal_words[250] = 32'b10001001010011011111001111001111;
        normal_words[251] = 32'b11010010011110001101110110111110;
        normal_words[252] = 32'b11111000011011110100001010100001;
        normal_words[253] = 32'b10001110000000000011001000110110;
        normal_words[254] = 32'b01101100000011001011110101000000;
        normal_words[255] = 32'b01000011011011101100011101000110;
        normal_words[256] = 32'b01101001001100111110010111010111;
        normal_words[257] = 32'b10100001000011110011101101100011;
        normal_words[258] = 32'b00110110100000100000110000100111;
        normal_words[259] = 32'b01011000111001100011110011110110;
        normal_words[260] = 32'b01000010110010011100001111110111;
        normal_words[261] = 32'b00010011111000001001101000101110;
        normal_words[262] = 32'b00101010100101011000000101110101;
        normal_words[263] = 32'b10011011011101000011000001100111;
        normal_words[264] = 32'b00000000111110001011000100110000;
        normal_words[265] = 32'b01001011100011011111100011010110;
        normal_words[266] = 32'b00011101011110100111011100001110;
        normal_words[267] = 32'b11110000001000001100011110010100;
        normal_words[268] = 32'b01000011110111001100011011111010;
        normal_words[269] = 32'b01100100011000000000010000010111;
        normal_words[270] = 32'b01101100111010010000001100000010;
        normal_words[271] = 32'b11111101111101010101010011101011;
        normal_words[272] = 32'b10010010111111111101001101011101;
        normal_words[273] = 32'b10010011110110110111111001111100;
        normal_words[274] = 32'b00111110111011101100011110111101;
        normal_words[275] = 32'b10000001000110011111011001010111;
        normal_words[276] = 32'b01010101011011101010011101111000;
        normal_words[277] = 32'b10100011011101011100101000110101;
        normal_words[278] = 32'b11001010010111010110010001100010;
        normal_words[279] = 32'b00101100000000110011101000110101;
        normal_words[280] = 32'b11110111011010100011000111100100;
        normal_words[281] = 32'b11011110100000011000100010100110;
        normal_words[282] = 32'b11000101001111101110010000100011;
        normal_words[283] = 32'b01011011110100111000110000111011;
        normal_words[284] = 32'b11001000101101010100010111111101;
        normal_words[285] = 32'b00001111100010011101100000001111;
        normal_words[286] = 32'b01001110000010100001100001000001;
        normal_words[287] = 32'b11111010111000010100001110101010;
        normal_words[288] = 32'b00111000100001111101101100100101;
        normal_words[289] = 32'b01101010100011111111010001110001;
        normal_words[290] = 32'b11111000010100110010011010000001;
        normal_words[291] = 32'b10111010011111000001010000110010;
        normal_words[292] = 32'b00110000101001110111000110011111;
        normal_words[293] = 32'b11001011111111010001010111000010;
        normal_words[294] = 32'b01110011000011010101110000000100;
        normal_words[295] = 32'b01100000011000100011111110100110;
        normal_words[296] = 32'b11001001100011111111000110100111;
        normal_words[297] = 32'b01111000111101001101010100010001;
        normal_words[298] = 32'b01110101100011010101011000110000;
        normal_words[299] = 32'b11010100000100001010101010111111;
        normal_words[300] = 32'b01011011100010011110101100000011;
        normal_words[301] = 32'b10101100011000001001111001111010;
        normal_words[302] = 32'b11011101010001000011101011110000;
        normal_words[303] = 32'b01101100000000001110100001011100;
        normal_words[304] = 32'b10000101011001100010000010001100;
        normal_words[305] = 32'b10100110100100110100001000100101;
        normal_words[306] = 32'b11101000100111100100010001010101;
        normal_words[307] = 32'b01010101101100111111000100111101;
        normal_words[308] = 32'b00101110110010111100111010011010;
        normal_words[309] = 32'b10010100101110100110101010000011;
        normal_words[310] = 32'b01101000011110000001010100110111;
        normal_words[311] = 32'b01000101110100100110100111011011;
        normal_words[312] = 32'b10001010000000001000110110001011;
        normal_words[313] = 32'b10111010001100111001011010101111;
        normal_words[314] = 32'b01011011110010100101110000011001;
        normal_words[315] = 32'b11011010101101011101101010000111;
        normal_words[316] = 32'b01110011100110111001011001111101;
        normal_words[317] = 32'b00010001100010101110010011101010;
        normal_words[318] = 32'b01001011000110111011111010000100;
        normal_words[319] = 32'b10101001101110000011010011110010;
        normal_words[320] = 32'b01000011101000001101000111010000;
        normal_words[321] = 32'b00100101001110100110000001100000;
        normal_words[322] = 32'b00101100111111111101110011110110;
        normal_words[323] = 32'b00110011000011001110001100100110;
        normal_words[324] = 32'b01100101001010000111001011001010;
        normal_words[325] = 32'b01011110010100100000101010010010;
        normal_words[326] = 32'b10011101110001011100110000100101;
        normal_words[327] = 32'b10000110110101000110111010011000;
        normal_words[328] = 32'b00000010100100111110001100111101;
        normal_words[329] = 32'b10111101110010010101000000111001;
        normal_words[330] = 32'b00101010011000010011011110110010;
        normal_words[331] = 32'b11111101011100110001101101100001;
        normal_words[332] = 32'b10001111111111001011101100111000;
        normal_words[333] = 32'b01000111011011011110001001111111;
        normal_words[334] = 32'b00100000000101000011101000110001;
        normal_words[335] = 32'b00000100100011000001100001111110;
        normal_words[336] = 32'b00001101110111100111000100100010;
        normal_words[337] = 32'b11101001100010110111101110010110;
        normal_words[338] = 32'b01011100011011111000010011110100;
        normal_words[339] = 32'b00010110111000001001011010010111;
        normal_words[340] = 32'b11000000100001010001100111101110;
        normal_words[341] = 32'b11111011111111101010110011110011;
        normal_words[342] = 32'b11000010011000110101111011000011;
        normal_words[343] = 32'b11100010100011011001101001011101;
        normal_words[344] = 32'b10110001011001111101110110110110;
        normal_words[345] = 32'b11100101100101001000111001010000;
        normal_words[346] = 32'b11110100110100000001101100011110;
        normal_words[347] = 32'b00010011110001001110011101010100;
        normal_words[348] = 32'b10010010101000011110000110010111;
        normal_words[349] = 32'b01000111001111100001101101111010;
        normal_words[350] = 32'b00101101111111001000001110101110;
        normal_words[351] = 32'b11010110001110110010110010000101;
        normal_words[352] = 32'b00101100000100110100000110010010;
        normal_words[353] = 32'b00100111100111101010011101001000;
        normal_words[354] = 32'b01001011000010010000101001001101;
        normal_words[355] = 32'b01111001110100100111010000101011;
        normal_words[356] = 32'b00010011000011110101011000100100;
        normal_words[357] = 32'b11000011110110101011010111011110;
        normal_words[358] = 32'b10011010111111000010111001111001;
        normal_words[359] = 32'b01111000000111010011111001001110;
        normal_words[360] = 32'b01001011001000011111011110010001;
        normal_words[361] = 32'b10111111010011000101010011010101;
        normal_words[362] = 32'b11001111000000110001000010100101;
        normal_words[363] = 32'b10010111101100100011001101100011;
        normal_words[364] = 32'b10011000000101001111001001100100;
        normal_words[365] = 32'b01001010110101000000010110001101;
        normal_words[366] = 32'b01010111010101100011101010101001;
        normal_words[367] = 32'b01100100101110000001010011110110;
        normal_words[368] = 32'b00100110100111100011011011111110;
        normal_words[369] = 32'b10110010101010001000010010110000;
        normal_words[370] = 32'b10100101111100110100111001101100;
        normal_words[371] = 32'b11011101001100101101011111110010;
        normal_words[372] = 32'b11010001011000011011001011101101;
        normal_words[373] = 32'b11111100001101001001110101000001;
        normal_words[374] = 32'b00001101100101010101111001111011;
        normal_words[375] = 32'b10011101010110011000101001101011;
        normal_words[376] = 32'b00100000110000100001111101100110;
        normal_words[377] = 32'b11010101101001110001010111010010;
        normal_words[378] = 32'b11000000100000111001001011001110;
        normal_words[379] = 32'b10110011111110100010010110001101;
        normal_words[380] = 32'b01110010001010101011001111101001;
        normal_words[381] = 32'b11000111011011011011101110111011;
        normal_words[382] = 32'b11000010010111111111111011110001;
        normal_words[383] = 32'b11110111011011011110011101000010;
        normal_words[384] = 32'b10100000100000111011111001100001;
        normal_words[385] = 32'b01110010011011011110100110001010;
        normal_words[386] = 32'b10100010100111000010101110110101;
        normal_words[387] = 32'b10100011001110110101101111100110;
        normal_words[388] = 32'b01000011111110000001011001111100;
        normal_words[389] = 32'b11111110011011110110111111110011;
        normal_words[390] = 32'b10110011000010010111111000010001;
        normal_words[391] = 32'b00110100001000011000000110000111;
        normal_words[392] = 32'b11000110100110010101010111000001;
        normal_words[393] = 32'b10011010110101000101100110111010;
        normal_words[394] = 32'b11100010011000001011000100100110;
        normal_words[395] = 32'b01001101011011011011111000101010;
        normal_words[396] = 32'b10000010000001110000100001000110;
        normal_words[397] = 32'b10101011000111110100110100110110;
        normal_words[398] = 32'b00100010101001110000000100010101;
        normal_words[399] = 32'b01011110000001000100010001110111;
        normal_words[400] = 32'b01011000011011010011010110000001;
        normal_words[401] = 32'b11001100101001010110001110010011;
        normal_words[402] = 32'b00111011101010001100101110011011;
        normal_words[403] = 32'b11111011010110110011100110000110;
        normal_words[404] = 32'b11111110111001111111000010001011;
        normal_words[405] = 32'b11100011111001000101000011010001;
        normal_words[406] = 32'b11001011111010000011011111110101;
        normal_words[407] = 32'b11101011100001111110111110010000;
        normal_words[408] = 32'b11100011111101001001101010001000;
        normal_words[409] = 32'b00111101001110101000100100000110;
        normal_words[410] = 32'b11010110010000111001110000000110;
        normal_words[411] = 32'b01011111111100111100100000110111;
        normal_words[412] = 32'b11001001110100010111010000111011;
        normal_words[413] = 32'b11100101000101100110000000001100;
        normal_words[414] = 32'b00111001100111111111101101010000;
        normal_words[415] = 32'b01110111000011001110111011010010;
        normal_words[416] = 32'b10001010001111011010000111110010;
        normal_words[417] = 32'b11000011011101111111101101110111;
        normal_words[418] = 32'b01001110100001010001100111000001;
        normal_words[419] = 32'b00110001010001100000010100000000;
        normal_words[420] = 32'b10000010110110000010000001011110;
        normal_words[421] = 32'b01010111111001001001001111110000;
        normal_words[422] = 32'b10011100001000010111000011100110;
        normal_words[423] = 32'b00100101101001101111011011000100;
        normal_words[424] = 32'b01110110111011001110101010110010;
        normal_words[425] = 32'b10100100100111001011001110110011;
        normal_words[426] = 32'b00001111101101011100101111000010;
        normal_words[427] = 32'b11110110100000101110110011110001;
        normal_words[428] = 32'b10101010111010111111001011000011;
        normal_words[429] = 32'b00100101110110010100000100001101;
        normal_words[430] = 32'b01001010000011000001011011110110;
        normal_words[431] = 32'b10111101010011011010111100100110;
        normal_words[432] = 32'b00100000010011010100101010101001;
        normal_words[433] = 32'b00000000101000111101101001000000;
        normal_words[434] = 32'b01100001000000001100110110101111;
        normal_words[435] = 32'b01101100100010101010111010000111;
        normal_words[436] = 32'b01101011010011101011110011101001;
        normal_words[437] = 32'b10011101111000111010111101011100;
        normal_words[438] = 32'b00011100100001010001101001111011;
        normal_words[439] = 32'b11111100010001100010010010101100;
        normal_words[440] = 32'b00001101000010011101110100011101;
        normal_words[441] = 32'b11111010001001001010100011101001;
        normal_words[442] = 32'b10000010000100110110001100001011;
        normal_words[443] = 32'b00100001000010100011110001011000;
        normal_words[444] = 32'b01100110101010001010000100111101;
        normal_words[445] = 32'b10001101101010101100101001101001;
        normal_words[446] = 32'b10010101010010010110011000101000;
        normal_words[447] = 32'b00001010110001110011100011111011;
        normal_words[448] = 32'b10010100100111100001010011001010;
        normal_words[449] = 32'b00100110010011110001001011111101;
        normal_words[450] = 32'b00101100001011110001010000111111;
        normal_words[451] = 32'b10011010000000110001000010010111;
        normal_words[452] = 32'b01001000001100101100010111100101;
        normal_words[453] = 32'b11101101101111101110111000110110;
        normal_words[454] = 32'b00110000111010101010010110111001;
        normal_words[455] = 32'b00111011110110000111010101111100;
        normal_words[456] = 32'b01101101010101101111010100101001;
        normal_words[457] = 32'b00000011000111100101000110010111;
        normal_words[458] = 32'b10101010111001000101100100101110;
        normal_words[459] = 32'b11010001101100000111010101010111;
        normal_words[460] = 32'b01100110010110011110110110000110;
        normal_words[461] = 32'b00110010010110000001001111110100;
        normal_words[462] = 32'b01011111011010001100100110101101;
        normal_words[463] = 32'b11111110011011100001010000001110;
        normal_words[464] = 32'b00011001111001101001001110110010;
        normal_words[465] = 32'b11000111000000111100001011111101;
        normal_words[466] = 32'b01101100000101010100100101111010;
        normal_words[467] = 32'b01100101111111111000010101001000;
        normal_words[468] = 32'b01111011001111001110101101001011;
        normal_words[469] = 32'b00001110100111010000100110111010;
        normal_words[470] = 32'b11011111011001110010000000101111;
        normal_words[471] = 32'b00001101010011010001100000000010;
        normal_words[472] = 32'b00110000100001010011111010001110;
        normal_words[473] = 32'b01111010000010010110111111100101;
        normal_words[474] = 32'b00101100001011010011110111111000;
        normal_words[475] = 32'b10110110010001000110111001100111;
        normal_words[476] = 32'b10001001101000011111010101100011;
        normal_words[477] = 32'b00101100111001010011000101001101;
        normal_words[478] = 32'b10010001110100101001101100110111;
        normal_words[479] = 32'b01110011001001101101101010101001;
        normal_words[480] = 32'b11101111110101100111000011101100;
        normal_words[481] = 32'b00001001110000000110101110011111;
        normal_words[482] = 32'b10000001011001101000100010011001;
        normal_words[483] = 32'b00010011000111011110100010110010;
        normal_words[484] = 32'b10100100011110000010000000001010;
        normal_words[485] = 32'b00011010001001110011011000110100;
        normal_words[486] = 32'b11110110001010010111001101000110;
        normal_words[487] = 32'b11000000000100110001111000000001;
        normal_words[488] = 32'b10010000010111100100101011000011;
        normal_words[489] = 32'b10110000100010101010110110111110;
        normal_words[490] = 32'b11001000010000111011110010101001;
        normal_words[491] = 32'b10101001100001011110100100000110;
        normal_words[492] = 32'b00110110100010010100101010011100;
        normal_words[493] = 32'b11100110111000000100011000010001;
        normal_words[494] = 32'b10000110011111100110011110111100;
        normal_words[495] = 32'b01010101011000000110001101001011;
        normal_words[496] = 32'b11010011111001011011110110010001;
        normal_words[497] = 32'b11100010001111010100001110000110;
        normal_words[498] = 32'b01110111000100100101111001011111;
        normal_words[499] = 32'b01011101000100100001111000101010;
        normal_words[500] = 32'b01100011000110010000001010100100;
        normal_words[501] = 32'b11010111001001001000111010111010;
        normal_words[502] = 32'b01010100010000100101000111011101;
        normal_words[503] = 32'b00011110111100011000001000010110;
        normal_words[504] = 32'b00100101111011111110110101100100;
        normal_words[505] = 32'b00111100000110010010111000101000;
        normal_words[506] = 32'b00000011011111110010001100110000;
        normal_words[507] = 32'b10110010100000110000010010111100;
        normal_words[508] = 32'b10100000000110011101000000011011;
        normal_words[509] = 32'b00011011111110110011110000110111;
        normal_words[510] = 32'b00101101001010100010011011001110;
        normal_words[511] = 32'b11011101000101000111001101100101;
        normal_words[512] = 32'b10110101110110110100111110011111;
        normal_words[513] = 32'b11011010011000110001100001110110;
        normal_words[514] = 32'b01101010001000101101000011111111;
        normal_words[515] = 32'b01111011010000110000110001101100;
        normal_words[516] = 32'b01100101100110011010100101010011;
        normal_words[517] = 32'b10010110101111111100010111111010;
        normal_words[518] = 32'b00001001000101001100110101000010;
        normal_words[519] = 32'b01000011000100001000101100011001;
        normal_words[520] = 32'b11110100011011101000000101010100;
        normal_words[521] = 32'b01000111000000001011101110000110;
        normal_words[522] = 32'b01110010100010011110011010010011;
        normal_words[523] = 32'b11100100010100101000010111100111;
        normal_words[524] = 32'b00100001111011111100100111001000;
        normal_words[525] = 32'b11110111101010100101101011100001;
        normal_words[526] = 32'b01001010001110000110000011101111;
        normal_words[527] = 32'b10101110000101000001110111101111;
        normal_words[528] = 32'b11110111110010101010001110110111;
        normal_words[529] = 32'b10111100000110100111010011011110;
        normal_words[530] = 32'b11011001010011001011011001100011;
        normal_words[531] = 32'b10010101011111101011111111000011;
        normal_words[532] = 32'b11000110110011100000111000101011;
        normal_words[533] = 32'b10001111010000110001000110011010;
        normal_words[534] = 32'b00000011000101000011001010000001;
        normal_words[535] = 32'b00001011100111101101010100110001;
        normal_words[536] = 32'b11101001010011011100111001110100;
        normal_words[537] = 32'b11000011011001011111111000101001;
        normal_words[538] = 32'b11100010011001000001010110100100;
        normal_words[539] = 32'b10011111010111100101010101001000;
        normal_words[540] = 32'b11111110011010101101010111101111;
        normal_words[541] = 32'b01000011001001001001100011111011;
        normal_words[542] = 32'b11001000101101111010010010100011;
        normal_words[543] = 32'b11110101111010110000011100011011;
        normal_words[544] = 32'b01101111011101110111010110111101;
        normal_words[545] = 32'b11110110001111010100011110100001;
        normal_words[546] = 32'b00111011010000101100001101000000;
        normal_words[547] = 32'b01010000100010000010110011111001;
        normal_words[548] = 32'b10010011011111010010111110100000;
        normal_words[549] = 32'b11110001000011000111101010110111;
        normal_words[550] = 32'b00110000111010101000111010001101;
        normal_words[551] = 32'b00010010011010110010010111010001;
        normal_words[552] = 32'b00000000000000000000000000010101;
        // Example bit positions from CSV (replace with actual data)

        // Initialize sparse pairs
        sparse_pairs[0] = {16'd148, 16'd342};
        sparse_pairs[1] = {16'd414, 16'd605};
        sparse_pairs[2] = {16'd627, 16'd1031};
        sparse_pairs[3] = {16'd1031, 16'd1435};
        sparse_pairs[4] = {16'd1478, 16'd1545};
        sparse_pairs[5] = {16'd1957, 16'd2201};
        sparse_pairs[6] = {16'd2201, 16'd2446};
        sparse_pairs[7] = {16'd2624, 16'd2794};
        sparse_pairs[8] = {16'd2794, 16'd2964};
        sparse_pairs[9] = {16'd3004, 16'd3015};
        sparse_pairs[10] = {16'd3037, 16'd3399};
        sparse_pairs[11] = {16'd3399, 16'd3761};
        sparse_pairs[12] = {16'd3761, 16'd4123};
        sparse_pairs[13] = {16'd4137, 16'd4166};
        sparse_pairs[14] = {16'd4167, 16'd4366};
        sparse_pairs[15] = {16'd4556, 16'd4690};
        sparse_pairs[16] = {16'd4690, 16'd4825};
        sparse_pairs[17] = {16'd6724, 16'd6816};
        sparse_pairs[18] = {16'd6913, 16'd7064};
        sparse_pairs[19] = {16'd7337, 16'd7526};
        sparse_pairs[20] = {16'd7848, 16'd8013};
        sparse_pairs[21] = {16'd8013, 16'd8179};
        sparse_pairs[22] = {16'd8463, 16'd8606};
        sparse_pairs[23] = {16'd8927, 16'd9048};
        sparse_pairs[24] = {16'd9048, 16'd9169};
        sparse_pairs[25] = {16'd9242, 16'd9552};
        sparse_pairs[26] = {16'd9552, 16'd9863};
        sparse_pairs[27] = {16'd9921, 16'd9924};
        sparse_pairs[28] = {16'd10272, 16'd10406};
        sparse_pairs[29] = {16'd10406, 16'd10540};
        sparse_pairs[30] = {16'd10560, 16'd10646};
        sparse_pairs[31] = {16'd10914, 16'd11115};
        sparse_pairs[32] = {16'd11115, 16'd11317};
        sparse_pairs[33] = {16'd11348, 16'd11458};
        sparse_pairs[34] = {16'd11458, 16'd11569};
        sparse_pairs[35] = {16'd12390, 16'd12640};
        sparse_pairs[36] = {16'd12640, 16'd12891};
        sparse_pairs[37] = {16'd13089, 16'd13117};
        sparse_pairs[38] = {16'd13120, 16'd13348};
        sparse_pairs[39] = {16'd13348, 16'd13577};
        sparse_pairs[40] = {16'd14633, 16'd14653};
        sparse_pairs[41] = {16'd14772, 16'd15122};
        sparse_pairs[42] = {16'd15122, 16'd15473};
        sparse_pairs[43] = {16'd15607, 16'd15690};
        sparse_pairs[44] = {16'd15761, 16'd15803};
        sparse_pairs[45] = {16'd16003, 16'd16262};
        sparse_pairs[46] = {16'd16262, 16'd16522};
        sparse_pairs[47] = {16'd16575, 16'd16721};
        sparse_pairs[48] = {16'd16721, 16'd16868};
        sparse_pairs[49] = {16'd16888, 16'd17336};
                
        rst_n = 0;
        start_process = 0;
        #(CLK_PERIOD * 2);
        rst_n = 1;
        #(CLK_PERIOD);


        for(pair_idx = 0; pair_idx < MEM_SPARSE_SIZE; pair_idx = pair_idx + 1) begin

            sparse_mem_addr_i = pair_idx;
            sparse_mem_data_i = sparse_pairs[pair_idx];
            start_process = 1;
            #(CLK_PERIOD);

            // Provide normal memory data when requested
            wait(normal_mem_addr_o == 0);
            #(CLK_PERIOD);
            normal_mem_data_i = normal_words[0];
            

            wait(normal_mem_addr_o == 551);
            #(CLK_PERIOD);
            normal_mem_data_i = normal_words[551];
                    

            wait(normal_mem_addr_o == 552);
            #(CLK_PERIOD);
            normal_mem_data_i = normal_words[552];
            
            

            acc_start_idx_high = sparse_mem_data_i[31:16] >> 5;  // 상위 16비트를 선택하고 32로 나눔
            acc_start_idx_low = sparse_mem_data_i[15:0] >> 5;    // 하위 16비트를 선택하고 32로 나눔

            high_low_diff = acc_start_idx_low - acc_start_idx_high;

            // Provide accumulator memory data based on acc_mem_addr_o
            wait(acc_mem_addr_o == acc_start_idx_high); // Wait for high shift address
            acc_mem_data_i = acc_words[acc_mem_addr_o]; // Initial acc data is 0
            
            #(CLK_PERIOD);
            
            
            wait(acc_mem_addr_o == acc_start_idx_low); // Wait for low shift address
            acc_mem_data_i = acc_words[acc_mem_addr_o]; // Initial acc data is 0
            
            #(CLK_PERIOD);
            

            #(CLK_PERIOD);



            // Wait for process_done signal before moving to next iteration
            wait(process_done);
            #(CLK_PERIOD * 2);
            rst_n = 0;
            start_process = 0;
            #(CLK_PERIOD * 2);
            rst_n = 1;
            #(CLK_PERIOD);
        end

        #(CLK_PERIOD);
        #(CLK_PERIOD);
        #(CLK_PERIOD);


        // Wait for process completion
        wait(process_done);
        #(CLK_PERIOD * 5);

        // Test completed
        $display("Test completed successfully!");
        $finish;
    end

    // Monitor acc_mem_write_en to update acc_words
    always @(posedge clk) begin
        if (acc_mem_write_en) begin
            acc_words[acc_mem_addr_o] <= acc_mem_write_data_o;
        end
    end

    // Monitor important signals
    initial begin
        $monitor("Time=%0t rst_n=%b start=%b busy=%b done=%b",
                 $time, rst_n, start_process, busy, process_done);
    end

endmodule