/* 
ChipWhisperer Artix Target - Simple testbench to check for signs of life.

Copyright (c) 2020, NewAE Technology Inc.
All rights reserved.

Redistribution and use in source and binary forms, with or without
modification, are permitted without restriction. Note that modules within
the project may have additional restrictions, please carefully inspect
additional licenses.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR
ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
(INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
(INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

The views and conclusions contained in the software and documentation are those
of the authors and should not be interpreted as representing official policies,
either expressed or implied, of NewAE Technology Inc.
*/

`timescale 1ns / 1ns
`default_nettype none 

`include "/home/boochoo/hqc/dummy-insertion-sparse-polymult/CW305/aes/cw305_aes_defines.v"

module tb();
    parameter pADDR_WIDTH = 21;
    parameter pBYTECNT_SIZE = 7;
    parameter pUSB_CLOCK_PERIOD = 10;
    parameter pPLL_CLOCK_PERIOD = 6;
    parameter pSEED = 1;
    parameter pTIMEOUT = 3000000;
    parameter pVERBOSE = 0;
    parameter pDUMP = 0;
    parameter WEIGHT = 2; //2
    parameter MEM_SIZE = 553;
   
    reg [32-1:0] normal_words [0:MEM_SIZE - 1];
    reg [15:0] sparse_pairs [0:WEIGHT-1];
    reg usb_clk;
    reg usb_clk_enable;
    wire [7:0] usb_data;
    reg [7:0] usb_wdata;
    reg [pADDR_WIDTH-1:0] usb_addr;
    reg usb_rdn;
    reg usb_wrn;
    reg usb_cen;
    reg usb_trigger;

    reg j16_sel;
    reg k16_sel;
    reg k15_sel;
    reg l14_sel;
    reg pushbutton;
    reg pll_clk1;
    wire tio_clkin;
    wire trig_out;

    wire led1;
    wire led2;
    wire led3;

    wire tio_trigger;
    wire tio_clkout;


    integer seed;
    integer errors;
    integer warnings;
    integer i;
    integer j;
    
    reg [31:0] write_data;

    wire clk = pll_clk1;  // shorthand for testbench

   integer cycle;
   integer total_time;

   reg [127:0] read_data;
   reg [127:0] expected_cipher = 128'h8a278bf8fa2812bc39e52c76205af377;

   reg [127:0] textin_extended;
   reg [127:0] key_extended;

   reg [127:0] textin_extended;
   reg [127:0] key_extended;

   task encrypt_index;
      input [15:0] textin;  // 16비트 입력값
      input [9:0] key;      // 8비트 정수 키 값
      begin

         // TEXTIN을 16비트에서 128비트로 확장 (상위 112비트는 0으로 패딩)
         textin_extended = {112'b0, textin};

         // KEY를 8비트 정수에서 128비트로 확장 (상위 120비트는 0으로 패딩)
         key_extended = {118'b0, key};

         // TEXTIN과 KEY를 레지스터에 저장
         write_bytes(0, 16, `REG_CRYPT_TEXTIN, textin_extended);
         write_bytes(0, 16, `REG_CRYPT_KEY, key_extended);

         $display("Encrypting via register...");
         write_byte(0, `REG_CRYPT_GO, 0, 1);
         repeat (5) @(posedge usb_clk);
         wait_done();
         read_bytes(0, 16, `REG_CRYPT_CIPHEROUT, read_data);

      end
   endtask

   task encrypt_text;
      input [31:0] textin;  // 16비트 입력값
      input [9:0] key;      // 8비트 정수 키 값
      begin

         // TEXTIN을 16비트에서 128비트로 확장 (상위 112비트는 0으로 패딩)
         textin_extended = {96'b0, textin};

         // KEY를 8비트 정수에서 128비트로 확장 (상위 120비트는 0으로 패딩)
         key_extended = {118'b0, key};

         // TEXTIN과 KEY를 레지스터에 저장
         write_bytes(0, 16, `REG_CRYPT_TEXTIN, textin_extended);
         write_bytes(0, 16, `REG_CRYPT_KEY, key_extended);

         $display("Encrypting via register...");
         write_byte(0, `REG_CRYPT_GO, 0, 1);
         repeat (5) @(posedge usb_clk);
         wait_done();
         read_bytes(0, 16, `REG_CRYPT_CIPHEROUT, read_data);

      end
   endtask


   task write_byte;
      input [1:0] block;
      input [pADDR_WIDTH-pBYTECNT_SIZE-1:0] address;
      input [pBYTECNT_SIZE-1:0] subbyte;
      input [7:0] data;
      begin
         @(posedge usb_clk);
         usb_addr = {block, address[5:0], subbyte};
         usb_wdata = data;
         usb_wrn = 0;
         @(posedge usb_clk);
         usb_cen = 0;
         @(posedge usb_clk);
         usb_cen = 1;
         @(posedge usb_clk);
         usb_wrn = 1;
         @(posedge usb_clk);
      end
   endtask


   task read_byte;
      input [1:0] block;
      input [pADDR_WIDTH-pBYTECNT_SIZE-1:0] address;
      input [pBYTECNT_SIZE-1:0] subbyte;
      output [7:0] data;
      begin
         @(posedge usb_clk);
         usb_addr = {block, address[5:0], subbyte};
         @(posedge usb_clk);
         usb_rdn = 0;
         usb_cen = 0;
         @(posedge usb_clk);
         @(posedge usb_clk);
         #1 data = usb_data;
         @(posedge usb_clk);
         usb_rdn = 1;
         usb_cen = 1;
         repeat(2) @(posedge usb_clk);
      end
   endtask


   task write_bytes;
      input [1:0] block;
      input [7:0] bytes;
      input [pADDR_WIDTH-pBYTECNT_SIZE-1:0] address;
      input [255:0] data;
      integer subbyte;
      begin
         for (subbyte = 0; subbyte < bytes; subbyte = subbyte + 1)
            write_byte(block, address, subbyte, data[subbyte*8 +: 8]);
         if (pVERBOSE)
            $display("Write %0h", data);
      end
   endtask


   task read_bytes;
      input [1:0] block;
      input [7:0] bytes;
      input [pADDR_WIDTH-pBYTECNT_SIZE-1:0] address;
      output [255:0] data;
      integer subbyte;
      begin
         for (subbyte = 0; subbyte < bytes; subbyte = subbyte + 1)
            read_byte(block, address, subbyte, data[subbyte*8 +: 8]);
         if (pVERBOSE)
            $display("Read %0h", data);
      end
   endtask




   initial begin


      normal_words[0] = 32'b01011110111001100110110110100101;
      normal_words[1] = 32'b01001011100010111011010011011000;
      normal_words[2] = 32'b11010000111001001101101101110100;
      normal_words[3] = 32'b11110100111010101100100010111111;
      normal_words[4] = 32'b10111111100011101100000110011100;
      normal_words[5] = 32'b00001100010010011101000111110101;
      normal_words[6] = 32'b00001000110001001010010000100110;
      normal_words[7] = 32'b10101011001011001010111001010010;
      normal_words[8] = 32'b00110111100100010010010110100010;
      normal_words[9] = 32'b11100110101010011111001101000111;
      normal_words[10] = 32'b11000111110100010001011001101100;
      normal_words[11] = 32'b11001001101100111100010000001000;
      normal_words[12] = 32'b10111010000000101011101100011011;
      normal_words[13] = 32'b11001011000111000110111010011111;
      normal_words[14] = 32'b10110111011100011001100011001110;
      normal_words[15] = 32'b10101011010101111101001100100001;
      normal_words[16] = 32'b01111001011101000001000100010110;
      normal_words[17] = 32'b10001100000100011010010010101010;
      normal_words[18] = 32'b00010100010010111001001010001001;
      normal_words[19] = 32'b01010111001000110000001100010010;
      normal_words[20] = 32'b10010000001111100100110000000100;
      normal_words[21] = 32'b00011010110110000000000000001100;
      normal_words[22] = 32'b01000111111111010000000000110010;
      normal_words[23] = 32'b01110010001100111101111101011001;
      normal_words[24] = 32'b10111110010000011010010100101000;
      normal_words[25] = 32'b00010011000010001000001011100000;
      normal_words[26] = 32'b00000111100001011010010011111000;
      normal_words[27] = 32'b10101001010001100000010010110101;
      normal_words[28] = 32'b11101010010111001101001111110111;
      normal_words[29] = 32'b11110111110011011011011111100001;
      normal_words[30] = 32'b11011101001000001010010000001011;
      normal_words[31] = 32'b01011000011011011100001101110100;
      normal_words[32] = 32'b11101010010011010101001110011000;
      normal_words[33] = 32'b10111000000111101110011001110011;
      normal_words[34] = 32'b11100100000101001010001010111100;
      normal_words[35] = 32'b01010100001110010110011000111100;
      normal_words[36] = 32'b01100101011100101111101101010000;
      normal_words[37] = 32'b10111101000110110000100001110001;
      normal_words[38] = 32'b01110111111111000010011010110010;
      normal_words[39] = 32'b01000000001011110111000010000100;
      normal_words[40] = 32'b10010000100000111001010110110101;
      normal_words[41] = 32'b11111110101011011100000000110100;
      normal_words[42] = 32'b00100011011010101110110101110111;
      normal_words[43] = 32'b01001111011011100100101110001101;
      normal_words[44] = 32'b10111100011110110101101011001001;
      normal_words[45] = 32'b11100011111010100010000100000001;
      normal_words[46] = 32'b10110111110101001111000101111000;
      normal_words[47] = 32'b01001011010001001100010010111001;
      normal_words[48] = 32'b01000110011001010011011101100101;
      normal_words[49] = 32'b01010111011000111101011101011011;
      normal_words[50] = 32'b11001000110100010101111110111001;
      normal_words[51] = 32'b01101111011010100001000111101001;
      normal_words[52] = 32'b10001110110100100111101110101111;
      normal_words[53] = 32'b10000110000000011011010001111000;
      normal_words[54] = 32'b10001000011111100110110100111110;
      normal_words[55] = 32'b01101100100100101001011111111111;
      normal_words[56] = 32'b00001100010111001001010100111101;
      normal_words[57] = 32'b11010111110111100101010110000000;
      normal_words[58] = 32'b00010011000011011001110111100011;
      normal_words[59] = 32'b01011111100001001101001001011000;
      normal_words[60] = 32'b01010110011110101000100000110110;
      normal_words[61] = 32'b01110010111100100001101001110100;
      normal_words[62] = 32'b01010100010011110110001010111011;
      normal_words[63] = 32'b10000011000111111011010001100011;
      normal_words[64] = 32'b10000111101101101011100100100111;
      normal_words[65] = 32'b01001100101000010010011110100110;
      normal_words[66] = 32'b11100101011100001101111001010101;
      normal_words[67] = 32'b11011100011011001100000100111001;
      normal_words[68] = 32'b10111000010000011000001010000100;
      normal_words[69] = 32'b11010010000000110010000101010111;
      normal_words[70] = 32'b01000000011100011110010010110101;
      normal_words[71] = 32'b00000000010001000100010100010011;
      normal_words[72] = 32'b00010010001110001111111011010100;
      normal_words[73] = 32'b10111100101000011001000010100001;
      normal_words[74] = 32'b00111111110110010011111110010010;
      normal_words[75] = 32'b10000010011010101110111011110110;
      normal_words[76] = 32'b01111000011001100011100011101111;
      normal_words[77] = 32'b01001010000001110001001011100011;
      normal_words[78] = 32'b10110010111111101110111010100100;
      normal_words[79] = 32'b00010011000100101110101000111011;
      normal_words[80] = 32'b11000100101011001101101100000111;
      normal_words[81] = 32'b11011101011110100101011001100111;
      normal_words[82] = 32'b10111010110111010000000110110011;
      normal_words[83] = 32'b11110011001110100001001001010000;
      normal_words[84] = 32'b11000101000000011100011011110011;
      normal_words[85] = 32'b11110001000100001010001001101000;
      normal_words[86] = 32'b01101101110000001100111111010001;
      normal_words[87] = 32'b10101000100011110010110101100111;
      normal_words[88] = 32'b11100110100011001111100010011111;
      normal_words[89] = 32'b01010011010000101110001011000000;
      normal_words[90] = 32'b11001011111000101001101111010100;
      normal_words[91] = 32'b01101011101001110001001010001110;
      normal_words[92] = 32'b10111110101101111010111111110110;
      normal_words[93] = 32'b00111111010100010010000101101011;
      normal_words[94] = 32'b10010111010001111111010111110110;
      normal_words[95] = 32'b00100001001101000100100101001010;
      normal_words[96] = 32'b01110001110011000011101000011000;
      normal_words[97] = 32'b01001101111111000110011110100110;
      normal_words[98] = 32'b10000011101110101010100000000011;
      normal_words[99] = 32'b01000000001101001100010100100110;
      normal_words[100] = 32'b01011111010100001001110000001000;
      normal_words[101] = 32'b01001010001001010111010000000011;
      normal_words[102] = 32'b10010010010100101100100111101100;
      normal_words[103] = 32'b10101101011000111111100011101100;
      normal_words[104] = 32'b11110000010011001110001111000110;
      normal_words[105] = 32'b00111111110010111000110010010011;
      normal_words[106] = 32'b00101010100011100111000111100000;
      normal_words[107] = 32'b01010101000000000000111101000000;
      normal_words[108] = 32'b00101111111000101101011011000101;
      normal_words[109] = 32'b10001100101111011010011000100111;
      normal_words[110] = 32'b00001010001111110101011110100011;
      normal_words[111] = 32'b11101000110010100110111001110111;
      normal_words[112] = 32'b11100001001111100110001001101010;
      normal_words[113] = 32'b00011011010100111011011100001000;
      normal_words[114] = 32'b10111000111110000100110110110100;
      normal_words[115] = 32'b00101100011100101100101001100010;
      normal_words[116] = 32'b11111001101101010001110110000010;
      normal_words[117] = 32'b01010010101101001101010010001111;
      normal_words[118] = 32'b00010110101110011111001101111000;
      normal_words[119] = 32'b01010100101011100000011110100001;
      normal_words[120] = 32'b11111001101100100010111100110110;
      normal_words[121] = 32'b01001010000111100101001011110011;
      normal_words[122] = 32'b01111010101010001000101010110110;
      normal_words[123] = 32'b11101100111011111100011001111100;
      normal_words[124] = 32'b10010011100001001010010101011101;
      normal_words[125] = 32'b11101001110000111110111110111000;
      normal_words[126] = 32'b10111000111111100110011000101001;
      normal_words[127] = 32'b00010000110001100000111110111011;
      normal_words[128] = 32'b10010011111001011101110001100011;
      normal_words[129] = 32'b11000000010001100000100110001101;
      normal_words[130] = 32'b01010101000101111011110011001100;
      normal_words[131] = 32'b01010110010011101111101010011101;
      normal_words[132] = 32'b10101101100101101000000011101001;
      normal_words[133] = 32'b11010001011110110000101100010010;
      normal_words[134] = 32'b01111100000000100110110000100111;
      normal_words[135] = 32'b01000100100100011011011011010001;
      normal_words[136] = 32'b11011110111111001100111100010011;
      normal_words[137] = 32'b10001101010000100011110000111001;
      normal_words[138] = 32'b00110110011011101100110110001011;
      normal_words[139] = 32'b10010010111001100100110001101101;
      normal_words[140] = 32'b10110001101011111101100100101111;
      normal_words[141] = 32'b00100011001100101011111000101111;
      normal_words[142] = 32'b00010101010010101000100110001110;
      normal_words[143] = 32'b01010001100110001001001010101001;
      normal_words[144] = 32'b10010000110000110110000000100101;
      normal_words[145] = 32'b11100100111001001111001110100011;
      normal_words[146] = 32'b00111110100110000000111000111110;
      normal_words[147] = 32'b10100001001100010110101100001111;
      normal_words[148] = 32'b01011010011100000110111001101001;
      normal_words[149] = 32'b11111100101100101101001110010101;
      normal_words[150] = 32'b11010111000111110100101101000101;
      normal_words[151] = 32'b00110101100001110110101000000110;
      normal_words[152] = 32'b00011000011111000011001011100011;
      normal_words[153] = 32'b10001100110111101111110101010101;
      normal_words[154] = 32'b10001101001100101110110111010111;
      normal_words[155] = 32'b11000010100011001111010111100011;
      normal_words[156] = 32'b00011000101111111110001010101111;
      normal_words[157] = 32'b10100101001101001000111111011000;
      normal_words[158] = 32'b10101100010100010101111011001001;
      normal_words[159] = 32'b00101110010110000100000110100000;
      normal_words[160] = 32'b10001000001011110000011100100001;
      normal_words[161] = 32'b00011110001001000001110000000001;
      normal_words[162] = 32'b10010010110100101011110001010110;
      normal_words[163] = 32'b01101010011000111100100101011100;
      normal_words[164] = 32'b00101010101110011101000111001101;
      normal_words[165] = 32'b10001111011001100101111110000100;
      normal_words[166] = 32'b11000010100011101110010000100111;
      normal_words[167] = 32'b00101011010000100110110011101010;
      normal_words[168] = 32'b10010110110100011111100111000111;
      normal_words[169] = 32'b10111001000111010000101011101101;
      normal_words[170] = 32'b10100101010100110110000000001110;
      normal_words[171] = 32'b00101001001011111100111011110111;
      normal_words[172] = 32'b11101110011110110001100011001100;
      normal_words[173] = 32'b01110010110000100111001000110111;
      normal_words[174] = 32'b01111001100101000000111010100001;
      normal_words[175] = 32'b01111010111111101101101000001001;
      normal_words[176] = 32'b00011100001110001000010111111001;
      normal_words[177] = 32'b11110011010011001110001101110100;
      normal_words[178] = 32'b00101000110000000110001100101100;
      normal_words[179] = 32'b00110010000100100111000000010111;
      normal_words[180] = 32'b11100001000101110001010110010111;
      normal_words[181] = 32'b01001010111100100011001001110110;
      normal_words[182] = 32'b11011100011110001101111010111111;
      normal_words[183] = 32'b01101100100001011101000000011111;
      normal_words[184] = 32'b00110010110011111000110110010010;
      normal_words[185] = 32'b00000000100100101100100100011001;
      normal_words[186] = 32'b10110000010011011101011001010101;
      normal_words[187] = 32'b01010110100000001100110010000000;
      normal_words[188] = 32'b00100111111010000011000110111010;
      normal_words[189] = 32'b11110101111010000111101111011000;
      normal_words[190] = 32'b10110110111111001111011111011000;
      normal_words[191] = 32'b10100010001011100100110110001111;
      normal_words[192] = 32'b00011011111111110001110010001010;
      normal_words[193] = 32'b10000001011001111101000000111010;
      normal_words[194] = 32'b00100110100000011011001011110110;
      normal_words[195] = 32'b00111000100111111110011011010101;
      normal_words[196] = 32'b01111111100100001011000111100011;
      normal_words[197] = 32'b11101000000100101010010000110111;
      normal_words[198] = 32'b01011110001000000001000000010111;
      normal_words[199] = 32'b11001100011110000000000010100011;
      normal_words[200] = 32'b01111100111101010111011110111100;
      normal_words[201] = 32'b11111011100000100111010100001001;
      normal_words[202] = 32'b01010111000011000100110000111111;
      normal_words[203] = 32'b10100101101000110011111001101001;
      normal_words[204] = 32'b10110011010011110101100011011010;
      normal_words[205] = 32'b11110111101101100000000101000010;
      normal_words[206] = 32'b01101100111101000001011011101100;
      normal_words[207] = 32'b00001001101010010000100000000100;
      normal_words[208] = 32'b01110111001000011010111001000110;
      normal_words[209] = 32'b00111000010110011010100101010001;
      normal_words[210] = 32'b11101110010000001110111000011110;
      normal_words[211] = 32'b10110011101101001010011010001001;
      normal_words[212] = 32'b01000100010101001110010011110001;
      normal_words[213] = 32'b00000010100111001000011100010100;
      normal_words[214] = 32'b00111000001010101101010001000000;
      normal_words[215] = 32'b11111011010101001100001100010101;
      normal_words[216] = 32'b01000100101110111010011100110100;
      normal_words[217] = 32'b10010100011111101010100001100110;
      normal_words[218] = 32'b11010000110111000010111000101101;
      normal_words[219] = 32'b11001001010000110101100010010100;
      normal_words[220] = 32'b01011101011110000001100110110000;
      normal_words[221] = 32'b10101001101001111101011010011101;
      normal_words[222] = 32'b10110010000101100011010111011011;
      normal_words[223] = 32'b00000011000110010101001100111111;
      normal_words[224] = 32'b10000001110111100001001101101000;
      normal_words[225] = 32'b01100100001001101111101110000011;
      normal_words[226] = 32'b01110001000000000011011111000100;
      normal_words[227] = 32'b00111111001010110010000100000011;
      normal_words[228] = 32'b00100100101100010101110001001101;
      normal_words[229] = 32'b11010110100010101111101001000101;
      normal_words[230] = 32'b00010100110101110011010110111000;
      normal_words[231] = 32'b10000001110101010001011111101100;
      normal_words[232] = 32'b00101110110001000010101000001010;
      normal_words[233] = 32'b01100001011011101010001101011111;
      normal_words[234] = 32'b11111011101101010111101001010010;
      normal_words[235] = 32'b01110010111010011100100110000101;
      normal_words[236] = 32'b00010100010101111011000101011111;
      normal_words[237] = 32'b10000001000000100101110000100101;
      normal_words[238] = 32'b01100010010100101111011101101111;
      normal_words[239] = 32'b00101110110000011010110000111010;
      normal_words[240] = 32'b00001100101011000101011111010110;
      normal_words[241] = 32'b00001011011110001010011111100000;
      normal_words[242] = 32'b01100110010011011011100011000001;
      normal_words[243] = 32'b01000000011011110011011101011011;
      normal_words[244] = 32'b01010011011010010000101010010100;
      normal_words[245] = 32'b10000110110101110110010011111100;
      normal_words[246] = 32'b11010001100110101010101001000000;
      normal_words[247] = 32'b11010010110010011000111000001100;
      normal_words[248] = 32'b01100000010101111101111101110111;
      normal_words[249] = 32'b11100000011110000111010011011111;
      normal_words[250] = 32'b11010111001110001011001111100001;
      normal_words[251] = 32'b11101000011100110101000011101000;
      normal_words[252] = 32'b00110000000100011001001100101000;
      normal_words[253] = 32'b00110000010000000011110101110101;
      normal_words[254] = 32'b11001000000111111011000110011010;
      normal_words[255] = 32'b01001101010111011010011101111001;
      normal_words[256] = 32'b11110111011011001010111000100010;
      normal_words[257] = 32'b11110101110010110001000001101110;
      normal_words[258] = 32'b10100100110011000000100001100000;
      normal_words[259] = 32'b00010010110010111010101001101011;
      normal_words[260] = 32'b00010001000011111000101011000011;
      normal_words[261] = 32'b00001000101101011111001101011111;
      normal_words[262] = 32'b11101110010110011001100101100000;
      normal_words[263] = 32'b10110110011110100011100011110100;
      normal_words[264] = 32'b10011010000010101000000101110111;
      normal_words[265] = 32'b00111111111111101100011110010011;
      normal_words[266] = 32'b11001000110110001110010101100010;
      normal_words[267] = 32'b01001100111010111100110000101101;
      normal_words[268] = 32'b10011001111100011100000000011001;
      normal_words[269] = 32'b11111000010011000010100100100011;
      normal_words[270] = 32'b10111010110010111111101101000000;
      normal_words[271] = 32'b00010011010101000101110110100010;
      normal_words[272] = 32'b01010000000111011011111011011011;
      normal_words[273] = 32'b10101110011011100111001010000000;
      normal_words[274] = 32'b11001001001101001101011000011001;
      normal_words[275] = 32'b00111101010100011100011100100111;
      normal_words[276] = 32'b11011101111110001001101011000011;
      normal_words[277] = 32'b01001100010010100010111101100110;
      normal_words[278] = 32'b00001110000100100111110110001010;
      normal_words[279] = 32'b10001001010111010001010001001000;
      normal_words[280] = 32'b01111101110011001000010001010010;
      normal_words[281] = 32'b00111101110101000101010000100000;
      normal_words[282] = 32'b01110010100111010000010100110011;
      normal_words[283] = 32'b01110001011111010011011100100110;
      normal_words[284] = 32'b10110010100011100011001110111100;
      normal_words[285] = 32'b11010001101110110011000110110100;
      normal_words[286] = 32'b10101001000111100001000000111111;
      normal_words[287] = 32'b01000111111100010101101111010100;
      normal_words[288] = 32'b00000110111011100010100011010110;
      normal_words[289] = 32'b00110011000111000011000010000011;
      normal_words[290] = 32'b00000111111010001111011111000011;
      normal_words[291] = 32'b10111011010101001001101111111111;
      normal_words[292] = 32'b11010111110101010000001001011000;
      normal_words[293] = 32'b10000101011000001011100101110101;
      normal_words[294] = 32'b10110110100010011100110011000111;
      normal_words[295] = 32'b10011010011010001101110011100001;
      normal_words[296] = 32'b10000111010110011111111101101000;
      normal_words[297] = 32'b10001100001010101111111110010101;
      normal_words[298] = 32'b10111011010001010001100101110010;
      normal_words[299] = 32'b10111101101110011101110011000000;
      normal_words[300] = 32'b00100111101010110101010100100101;
      normal_words[301] = 32'b11010101000110101010101101001100;
      normal_words[302] = 32'b10001111101001001010010110101001;
      normal_words[303] = 32'b11110111000010111010101101111011;
      normal_words[304] = 32'b10011001111100010100010110011011;
      normal_words[305] = 32'b01110100011010110001010110001110;
      normal_words[306] = 32'b00001101011011101110010001001111;
      normal_words[307] = 32'b11010111110110011000000101010111;
      normal_words[308] = 32'b01101000000001100001001101110110;
      normal_words[309] = 32'b11001100101011000101000110001010;
      normal_words[310] = 32'b10001100111001111000110010110111;
      normal_words[311] = 32'b00111010111111010001101101111110;
      normal_words[312] = 32'b10101000010100101100100110111101;
      normal_words[313] = 32'b00111000110100000100110011100100;
      normal_words[314] = 32'b10110000111010110101010001000011;
      normal_words[315] = 32'b11011110000110100000001100011000;
      normal_words[316] = 32'b01000001001001010010100100010000;
      normal_words[317] = 32'b10010101000101111000111101011010;
      normal_words[318] = 32'b10100011001100110011001111110000;
      normal_words[319] = 32'b00010101011001110010011101110101;
      normal_words[320] = 32'b00001010001000000100111111110000;
      normal_words[321] = 32'b01100101010111010000001001001010;
      normal_words[322] = 32'b00101101000111101001111100100000;
      normal_words[323] = 32'b01111111011110100010011100000111;
      normal_words[324] = 32'b11000100011111110010010001001111;
      normal_words[325] = 32'b11100100011001011110000110100011;
      normal_words[326] = 32'b10011110000101110011110101100011;
      normal_words[327] = 32'b11110111011101111011011000101111;
      normal_words[328] = 32'b01011010010010101000111111111000;
      normal_words[329] = 32'b10100101110101011111001011001100;
      normal_words[330] = 32'b11100011001100111110011000101100;
      normal_words[331] = 32'b11001111100100000101011010010110;
      normal_words[332] = 32'b00100001101100110101110100011000;
      normal_words[333] = 32'b01011100111011111000011100010101;
      normal_words[334] = 32'b11001101001111111000110100110010;
      normal_words[335] = 32'b10100100000001010110100010110110;
      normal_words[336] = 32'b00111111011100111010110010000010;
      normal_words[337] = 32'b00010101100010001100010000001110;
      normal_words[338] = 32'b01010001010011011111000001110101;
      normal_words[339] = 32'b10111101100100110000111011100000;
      normal_words[340] = 32'b00100000000101000011010100110011;
      normal_words[341] = 32'b10010000100010010011110011011100;
      normal_words[342] = 32'b00111111011000100100000010110000;
      normal_words[343] = 32'b11100100011100001010001111101010;
      normal_words[344] = 32'b10010001100111001111110010010111;
      normal_words[345] = 32'b11001010101000011101101001101000;
      normal_words[346] = 32'b01100110010000000011011100100000;
      normal_words[347] = 32'b01110111111101101000110001111111;
      normal_words[348] = 32'b11011011000110010111100000110101;
      normal_words[349] = 32'b00001101101010111011000010010100;
      normal_words[350] = 32'b01111001101101010101110101110001;
      normal_words[351] = 32'b00111001001100000101000011110100;
      normal_words[352] = 32'b11011110000011001001110011011101;
      normal_words[353] = 32'b10100110101111001100000110111101;
      normal_words[354] = 32'b01001001101101001111110101011101;
      normal_words[355] = 32'b00110011100100010111111111001001;
      normal_words[356] = 32'b11011110101100000111100110000010;
      normal_words[357] = 32'b01000000101101110111010000001100;
      normal_words[358] = 32'b10001001110111010011101011101000;
      normal_words[359] = 32'b10010111011000001101110001011001;
      normal_words[360] = 32'b01110011101111011110000110001101;
      normal_words[361] = 32'b11011101110011110000100110001000;
      normal_words[362] = 32'b10001010100101000111011100100010;
      normal_words[363] = 32'b01010101000101011111101101000101;
      normal_words[364] = 32'b01000011011101010001101001000001;
      normal_words[365] = 32'b01111100101110101001111111100111;
      normal_words[366] = 32'b11111011101000011110100010101010;
      normal_words[367] = 32'b01110010110101010101110110001001;
      normal_words[368] = 32'b11010000011111010001101100100011;
      normal_words[369] = 32'b11001111000000010100010010011110;
      normal_words[370] = 32'b10011100100111111110011100011111;
      normal_words[371] = 32'b00000100111001011000110110011110;
      normal_words[372] = 32'b10010101001101010110001011000111;
      normal_words[373] = 32'b11111010111110101000010010111100;
      normal_words[374] = 32'b11101111100100110010011010101101;
      normal_words[375] = 32'b01000011000100010001111010001100;
      normal_words[376] = 32'b00111001101010110010100100110111;
      normal_words[377] = 32'b11011000010010101010010011100111;
      normal_words[378] = 32'b00001100101111010110100010011110;
      normal_words[379] = 32'b00110000010101101101111101000000;
      normal_words[380] = 32'b10010100011000110111110010100000;
      normal_words[381] = 32'b00110111110101001101110111000001;
      normal_words[382] = 32'b11010101010000100101111010011000;
      normal_words[383] = 32'b01011110111111000110010101011010;
      normal_words[384] = 32'b10011100001100011011110110100100;
      normal_words[385] = 32'b11001011011010111111000110011010;
      normal_words[386] = 32'b10010001001100001011110011110010;
      normal_words[387] = 32'b10001001010001010010111111101001;
      normal_words[388] = 32'b01011100011111001110100000101100;
      normal_words[389] = 32'b00001011010001001011100101000000;
      normal_words[390] = 32'b11010110011010011000010010100000;
      normal_words[391] = 32'b01111111001111111011010100111010;
      normal_words[392] = 32'b11110101010011110111000000001111;
      normal_words[393] = 32'b11100011110100000001111100011011;
      normal_words[394] = 32'b11100000011001101000010000100000;
      normal_words[395] = 32'b10001011011010101111100001101011;
      normal_words[396] = 32'b00000111100100100110000100101000;
      normal_words[397] = 32'b01100111110011001010011101101101;
      normal_words[398] = 32'b10100110101001101001010010110001;
      normal_words[399] = 32'b00101000101101111011100111010000;
      normal_words[400] = 32'b01010100011000111101011111001101;
      normal_words[401] = 32'b00000111001010011000001101001101;
      normal_words[402] = 32'b01001101011000110011000001100100;
      normal_words[403] = 32'b01110000110101111111000111000110;
      normal_words[404] = 32'b00001010000100101011100101010011;
      normal_words[405] = 32'b11110111000011101011100011011000;
      normal_words[406] = 32'b11101000111111110011000010010101;
      normal_words[407] = 32'b10111111010111111100101100111100;
      normal_words[408] = 32'b00100011010010101101111101110001;
      normal_words[409] = 32'b00100011111010010001001000110101;
      normal_words[410] = 32'b11110101101100011111010100010111;
      normal_words[411] = 32'b11100000100101101100100101001010;
      normal_words[412] = 32'b01011011000001111110111100010100;
      normal_words[413] = 32'b01100111011110110000000101100001;
      normal_words[414] = 32'b10001000110011001111000001011000;
      normal_words[415] = 32'b11011000000000110101001010100011;
      normal_words[416] = 32'b11011100001111110010110011011111;
      normal_words[417] = 32'b11100101001000001100010101001100;
      normal_words[418] = 32'b01110110000100101101001101010101;
      normal_words[419] = 32'b11110110100011101000011111101101;
      normal_words[420] = 32'b01101000000000101101000101010100;
      normal_words[421] = 32'b01010010001000101101101001011001;
      normal_words[422] = 32'b00001111101011011101100001001100;
      normal_words[423] = 32'b00000001111000000011111011011111;
      normal_words[424] = 32'b11110011010010011101101001111010;
      normal_words[425] = 32'b00111000101000100010001011111101;
      normal_words[426] = 32'b11011011100000100100000110011011;
      normal_words[427] = 32'b01011011110111000101011111011100;
      normal_words[428] = 32'b10110001001100101010011110110000;
      normal_words[429] = 32'b10010001111111000110000101000011;
      normal_words[430] = 32'b11011101010010000010101000111110;
      normal_words[431] = 32'b10010101101001111101101110110001;
      normal_words[432] = 32'b00101011101101110100110110011011;
      normal_words[433] = 32'b10010100101010010011111101010100;
      normal_words[434] = 32'b11110011011000001101100101010001;
      normal_words[435] = 32'b01011111100110110010101100001011;
      normal_words[436] = 32'b10011111001111010000000000111100;
      normal_words[437] = 32'b10110010010110011000000101110110;
      normal_words[438] = 32'b10101011011011010100001010001110;
      normal_words[439] = 32'b11101110000100100000101001110000;
      normal_words[440] = 32'b10001001001110111101011010000010;
      normal_words[441] = 32'b10100110110001011001110110001011;
      normal_words[442] = 32'b00100111010001001000010011001001;
      normal_words[443] = 32'b01110111011101110100011110010110;
      normal_words[444] = 32'b10001101010101111100001000110011;
      normal_words[445] = 32'b10000011010000111101011111110010;
      normal_words[446] = 32'b10101011110011110001001101111110;
      normal_words[447] = 32'b11000110000011100011111110011011;
      normal_words[448] = 32'b10011111000110001100001000110100;
      normal_words[449] = 32'b11000010101000000111111111000110;
      normal_words[450] = 32'b00100001011010100011100100100101;
      normal_words[451] = 32'b11011111110000100011010111011000;
      normal_words[452] = 32'b10011100111001010111000111100000;
      normal_words[453] = 32'b01101100000000001111011001000110;
      normal_words[454] = 32'b10001101101001100011101111110001;
      normal_words[455] = 32'b01101011111001000010110111111100;
      normal_words[456] = 32'b10110100101011000010000110010010;
      normal_words[457] = 32'b01011101100110110010111110001100;
      normal_words[458] = 32'b10100101010110111110101001010111;
      normal_words[459] = 32'b11001101010011111010001111101111;
      normal_words[460] = 32'b10101000011011110001110111110111;
      normal_words[461] = 32'b11010110111111111111011101011010;
      normal_words[462] = 32'b01001110100000010000100010011000;
      normal_words[463] = 32'b00010010111010110010010100000100;
      normal_words[464] = 32'b11000110010101000000010111100111;
      normal_words[465] = 32'b10101000001010111011001000110011;
      normal_words[466] = 32'b00011111110101101000101001100100;
      normal_words[467] = 32'b01100001100100101000101101000110;
      normal_words[468] = 32'b00101000000101001001010001000100;
      normal_words[469] = 32'b10111110110110101011011101100100;
      normal_words[470] = 32'b00001011100110111110011010110110;
      normal_words[471] = 32'b00001011001001101001010001011001;
      normal_words[472] = 32'b11010000110100100010110001001101;
      normal_words[473] = 32'b01000100000111110101011001110001;
      normal_words[474] = 32'b00010001011010001001010110001111;
      normal_words[475] = 32'b11000011010010011101100100110111;
      normal_words[476] = 32'b10110001001001000001111100001010;
      normal_words[477] = 32'b11001010011011000001110001110011;
      normal_words[478] = 32'b11100011001100110000100010011000;
      normal_words[479] = 32'b01000001001100010100100001011000;
      normal_words[480] = 32'b01001011110001010000001010000000;
      normal_words[481] = 32'b01001011101011101001000100110100;
      normal_words[482] = 32'b00001000110000010101011001111001;
      normal_words[483] = 32'b10100011011110011111100101001011;
      normal_words[484] = 32'b01001001001100010000011111101001;
      normal_words[485] = 32'b11100100001001001000001011000010;
      normal_words[486] = 32'b10011111011010111101100001100011;
      normal_words[487] = 32'b10100101001001001100101010110100;
      normal_words[488] = 32'b11000001001111100011000101101101;
      normal_words[489] = 32'b00101101011101011100001000100000;
      normal_words[490] = 32'b11111010000000110000010100010111;
      normal_words[491] = 32'b11111110111110011110010111100010;
      normal_words[492] = 32'b11110100000111101100000111100010;
      normal_words[493] = 32'b10110000011011111010001101010000;
      normal_words[494] = 32'b00010001000000001110101111001101;
      normal_words[495] = 32'b10001001010111101100001110100000;
      normal_words[496] = 32'b11110101011100000111011001011110;
      normal_words[497] = 32'b01001010111100010001001101100010;
      normal_words[498] = 32'b01010001010101100101011110000100;
      normal_words[499] = 32'b11011100101000000000011100100100;
      normal_words[500] = 32'b11000010001001111001011000101001;
      normal_words[501] = 32'b10110100010111010000001111000110;
      normal_words[502] = 32'b01010001011101000001010111101011;
      normal_words[503] = 32'b10000011110011100101100001110001;
      normal_words[504] = 32'b00101110100110101100101111000010;
      normal_words[505] = 32'b10101010000110110011111000000110;
      normal_words[506] = 32'b00010010000110011011110010101010;
      normal_words[507] = 32'b01010011000011101111111010011101;
      normal_words[508] = 32'b11000110001101110111011101101101;
      normal_words[509] = 32'b00101110011111010110000110000100;
      normal_words[510] = 32'b01100010101110010011001100010010;
      normal_words[511] = 32'b00001100110010011101101111111100;
      normal_words[512] = 32'b11000101101110110010001100100100;
      normal_words[513] = 32'b11110100011011111001010101010111;
      normal_words[514] = 32'b01110101101111100110110010100010;
      normal_words[515] = 32'b01011100111001101011110100101110;
      normal_words[516] = 32'b00110010110101010001000110001110;
      normal_words[517] = 32'b11110111110111000100001000011101;
      normal_words[518] = 32'b00001010110101100001011101010010;
      normal_words[519] = 32'b10101111101111010010000111001011;
      normal_words[520] = 32'b10011010000000011001101110110101;
      normal_words[521] = 32'b00001001110110111100001111100000;
      normal_words[522] = 32'b10111101000011110011000100001100;
      normal_words[523] = 32'b11100011010010000001110101001000;
      normal_words[524] = 32'b00010101101010011011011110001001;
      normal_words[525] = 32'b11110000110100101100111001011101;
      normal_words[526] = 32'b11110111111010010010000011011011;
      normal_words[527] = 32'b11011011111111011111010110011001;
      normal_words[528] = 32'b10100100010110110100101100000110;
      normal_words[529] = 32'b00100010001010011101001111000001;
      normal_words[530] = 32'b10101111101001010111110011000000;
      normal_words[531] = 32'b10011100110100000010010011100000;
      normal_words[532] = 32'b11110100001001111010110011001000;
      normal_words[533] = 32'b01011100010011011100110010011010;
      normal_words[534] = 32'b01000011100000100000010011010110;
      normal_words[535] = 32'b10011001100101001101110001111111;
      normal_words[536] = 32'b01011101111010010110000010111001;
      normal_words[537] = 32'b01100100100111100111111111010111;
      normal_words[538] = 32'b01100001101100101001100100101101;
      normal_words[539] = 32'b01011111111011011000001000011111;
      normal_words[540] = 32'b11100110000101110000101110000000;
      normal_words[541] = 32'b01011001100000111001001011101100;
      normal_words[542] = 32'b00010000110111010111001100011111;
      normal_words[543] = 32'b01000011110001000110111000110100;
      normal_words[544] = 32'b00011111010001110000000010100011;
      normal_words[545] = 32'b10000010000010001000011110000001;
      normal_words[546] = 32'b00111101010011110101111010001000;
      normal_words[547] = 32'b01001001111100000011011111001011;
      normal_words[548] = 32'b01111110001101011111011111110100;
      normal_words[549] = 32'b01110100001001011010111001001010;
      normal_words[550] = 32'b01011111000110001011111111101111;
      normal_words[551] = 32'b01011101000001101000010001000100;
      normal_words[552] = 32'b00000000000000000000000000011110;

      sparse_pairs[0]  = 16'b0000000010010100;
      sparse_pairs[1]  = 16'b0000000101010110;
      sparse_pairs[2]  = 16'b0000000110011110;
      sparse_pairs[3]  = 16'b0000001001011101;
      sparse_pairs[4]  = 16'b0000001001110011;
      sparse_pairs[5]  = 16'b0000010110011011;
      sparse_pairs[6]  = 16'b0000010111000110;
      sparse_pairs[7]  = 16'b0000011000001001;
      sparse_pairs[8]  = 16'b0000011110100101;
      sparse_pairs[9]  = 16'b0000100110001110;
      sparse_pairs[10] = 16'b0000101001000000;
      sparse_pairs[11] = 16'b0000101110010100;
      sparse_pairs[12] = 16'b0000101110111100;
      sparse_pairs[13] = 16'b0000101111000111;
      sparse_pairs[14] = 16'b0000101111011101;
      sparse_pairs[15] = 16'b0001000000011011;
      sparse_pairs[16] = 16'b0001000000101001;
      sparse_pairs[17] = 16'b0001000001000110;
      sparse_pairs[18] = 16'b0001000001000111;
      sparse_pairs[19] = 16'b0001000100001110;
      sparse_pairs[20] = 16'b0001000111001100;
      sparse_pairs[21] = 16'b0001001011011001;
      sparse_pairs[22] = 16'b0001101001000100;
      sparse_pairs[23] = 16'b0001101010100000;
      sparse_pairs[24] = 16'b0001101100000001;
      sparse_pairs[25] = 16'b0001101110011000;
      sparse_pairs[26] = 16'b0001110010101001;
      sparse_pairs[27] = 16'b0001110101100110;
      sparse_pairs[28] = 16'b0001111010101000;
      sparse_pairs[29] = 16'b0001111111110011;
      sparse_pairs[30] = 16'b0010000100001111;
      sparse_pairs[31] = 16'b0010000110011110;
      sparse_pairs[32] = 16'b0010001011011111;
      sparse_pairs[33] = 16'b0010001111010001;
      sparse_pairs[34] = 16'b0010010000011010;
      sparse_pairs[35] = 16'b0010011010000111;
      sparse_pairs[36] = 16'b0010011011000001;
      sparse_pairs[37] = 16'b0010011011000100;
      sparse_pairs[38] = 16'b0010100000100000;
      sparse_pairs[39] = 16'b0010100100101100;
      sparse_pairs[40] = 16'b0010100101000000;
      sparse_pairs[41] = 16'b0010100110010110;
      sparse_pairs[42] = 16'b0010101010100010;
      sparse_pairs[43] = 16'b0010110000110101;
      sparse_pairs[44] = 16'b0010110001010100;
      sparse_pairs[45] = 16'b0010110100110001;
      sparse_pairs[46] = 16'b0011000001100110;
      sparse_pairs[47] = 16'b0011001001011011;
      sparse_pairs[48] = 16'b0011001100100001;
      sparse_pairs[49] = 16'b0011001100111101;
      sparse_pairs[50] = 16'b0011001101000000;
      sparse_pairs[51] = 16'b0011010100001001;
      sparse_pairs[52] = 16'b0011100100101001;
      sparse_pairs[53] = 16'b0011100100111101;
      sparse_pairs[54] = 16'b0011100110110100;
      sparse_pairs[55] = 16'b0011110001110001;
      sparse_pairs[56] = 16'b0011110011110111;
      sparse_pairs[57] = 16'b0011110101001010;
      sparse_pairs[58] = 16'b0011110110010001;
      sparse_pairs[59] = 16'b0011110110111011;
      sparse_pairs[60] = 16'b0011111010000011;
      sparse_pairs[61] = 16'b0100000010001010;
      sparse_pairs[62] = 16'b0100000010111111;
      sparse_pairs[63] = 16'b0100000111100100;
      sparse_pairs[64] = 16'b0100000111111000;
      sparse_pairs[65] = 16'b0100001110111000;


      // sparse_pairs[0]  = 16'b0000000001010100;
      // sparse_pairs[1]  = 16'b0000000011110101;
      // sparse_pairs[2]  = 16'b0000000100010010;
      // sparse_pairs[3]  = 16'b0000000110001010;
      // sparse_pairs[4]  = 16'b0000000111000010;
      // sparse_pairs[5]  = 16'b0000001001010101;
      // sparse_pairs[6]  = 16'b0000001101100100;
      // sparse_pairs[7]  = 16'b0000001111100101;
      // sparse_pairs[8]  = 16'b0000010001011000;
      // sparse_pairs[9]  = 16'b0000010101110000;
      // sparse_pairs[10] = 16'b0000010111111101;
      // sparse_pairs[11] = 16'b0000011000011110;
      // sparse_pairs[12] = 16'b0000011001101111;
      // sparse_pairs[13] = 16'b0000100101000100;
      // sparse_pairs[14] = 16'b0000101010001011;
      // sparse_pairs[15] = 16'b0000101111010010;
      // sparse_pairs[16] = 16'b0000101111101100;
      // sparse_pairs[17] = 16'b0000110001000010;
      // sparse_pairs[18] = 16'b0001000011010010;
      // sparse_pairs[19] = 16'b0001000101110010;
      // sparse_pairs[20] = 16'b0001000110000001;
      // sparse_pairs[21] = 16'b0001001000100001;
      // sparse_pairs[22] = 16'b0001001001010110;
      // sparse_pairs[23] = 16'b0001001010110111;
      // sparse_pairs[24] = 16'b0001001110010100;
      // sparse_pairs[25] = 16'b0001010001011100;
      // sparse_pairs[26] = 16'b0001010011100111;
      // sparse_pairs[27] = 16'b0001010111000011;
      // sparse_pairs[28] = 16'b0001011001000100;
      // sparse_pairs[29] = 16'b0010110110101001;
      // sparse_pairs[30] = 16'b0010111000010100;
      // sparse_pairs[31] = 16'b0010111011011110;
      // sparse_pairs[32] = 16'b0010111111001110;
      // sparse_pairs[33] = 16'b0011000011010010;
      // sparse_pairs[34] = 16'b0011000011010110;
      // sparse_pairs[35] = 16'b0011000100000110;
      // sparse_pairs[36] = 16'b0011001001010001;
      // sparse_pairs[37] = 16'b0011001100101011;
      // sparse_pairs[38] = 16'b0011001111001000;
      // sparse_pairs[39] = 16'b0011010011100011;
      // sparse_pairs[40] = 16'b0011010101100010;
      // sparse_pairs[41] = 16'b0011100010110100;
      // sparse_pairs[42] = 16'b0011100011101001;
      // sparse_pairs[43] = 16'b0011100100000110;
      // sparse_pairs[44] = 16'b0011100100111110;
      // sparse_pairs[45] = 16'b0011100111010010;
      // sparse_pairs[46] = 16'b0011101100001011;
      // sparse_pairs[47] = 16'b0011101101010011;
      // sparse_pairs[48] = 16'b0011101101101100;
      // sparse_pairs[49] = 16'b0011101111000101;
      // sparse_pairs[50] = 16'b0011110010010010;
      // sparse_pairs[51] = 16'b0011111000100001;
      // sparse_pairs[52] = 16'b0011111000101011;
      // sparse_pairs[53] = 16'b0011111100100101;
      // sparse_pairs[54] = 16'b0011111101101101;
      // sparse_pairs[55] = 16'b0100000001001110;
      // sparse_pairs[56] = 16'b0100000001001111;
      // sparse_pairs[57] = 16'b0100000101101011;
      // sparse_pairs[58] = 16'b0100000110111100;
      // sparse_pairs[59] = 16'b0100001000001010;
      // sparse_pairs[60] = 16'b0100001000110111;
      // sparse_pairs[61] = 16'b0100001010010000;
      // sparse_pairs[62] = 16'b0100001010010011;
      // sparse_pairs[63] = 16'b0100001110001001;
      // sparse_pairs[64] = 16'b0100010001000000;
      // sparse_pairs[65] = 16'b0100010011101000;

      seed = pSEED;
      errors = 0;
      warnings = 0;
      $display("Running with seed=%0d", seed);
      seed = $random;
      if (pDUMP) begin
         $dumpfile("results/tb.fst");
         $dumpvars(0, tb);
      end
      usb_clk = 1'b1;
      usb_clk_enable = 1'b1;
      pll_clk1 = 1'b1;

      usb_wdata = 0;
      usb_addr = 0;
      usb_rdn = 1;
      usb_wrn = 1;
      usb_cen = 1;
      usb_trigger = 0;

      j16_sel = 0;
      k16_sel = 0;
      k15_sel = 0;
      l14_sel = 0;
      pushbutton = 1;
      pll_clk1 = 0;

      #(pUSB_CLOCK_PERIOD*2) pushbutton = 0;
      #(pUSB_CLOCK_PERIOD*2) pushbutton = 1;
      #(pUSB_CLOCK_PERIOD*10);

      for (j = 0; j < WEIGHT; j = j + 1) begin
         encrypt_index(sparse_pairs[j], j);  // sparse_pairs[i]를 TEXTIN으로 사용, key 값은 i (0~65)
      end

      for (j =WEIGHT; j < MEM_SIZE + WEIGHT; j = j + 1) begin
         encrypt_text(normal_words[j - WEIGHT], j);  // normal_words[i-66]를 TEXTIN으로 사용, key 값은 i (66~618)
      end

      write_bytes(0, 16, `REG_CRYPT_TEXTIN, {32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF, 32'hFFFFFFFF});
      write_bytes(0, 16, `REG_CRYPT_KEY, {32'h80000000, 32'h0, 32'h0, 32'hFFFFFFFF});


      #(pUSB_CLOCK_PERIOD*2) pushbutton = 0;
      #(pUSB_CLOCK_PERIOD*2) pushbutton = 1;


      $display("Encrypting via register...");
      write_byte(0, `REG_CRYPT_GO, 0, 1);
      repeat (5) @(posedge usb_clk);
      wait_done();
      read_bytes(0, 16, `REG_CRYPT_CIPHEROUT, read_data);
      if (read_data == expected_cipher) begin
         $display("Good result");
      end
      else begin
         errors = errors + 1;
         $display("ERROR: expected %h", expected_cipher);
         $display("            got %h", read_data);
      end

      // normal_words[0] = 32'b01111000110101101010100101010101;
      // normal_words[1] = 32'b10100001101000110110101000010011;
      // normal_words[2] = 32'b11111011100000010110010101110001;
      // normal_words[3] = 32'b11010000111001110000010000100100;
      // normal_words[4] = 32'b01010101110110001111110010011010;
      // normal_words[5] = 32'b01011011000000011011001100111000;
      // normal_words[6] = 32'b10100001111111011100011111100100;
      // normal_words[7] = 32'b10111000111010001101010110101101;
      // normal_words[8] = 32'b00100111001000111111101101010000;
      // normal_words[9] = 32'b00010000010001011101010000111110;
      // normal_words[10] = 32'b11100100111010100111010001110000;
      // normal_words[11] = 32'b00010100011001010100101111111000;
      // normal_words[12] = 32'b00100011010110011001010011011101;
      // normal_words[13] = 32'b00100011001001010111011000001000;
      // normal_words[14] = 32'b10110100000111100001101100011000;
      // normal_words[15] = 32'b11010100101111101100100010001000;
      // normal_words[16] = 32'b01011001111100101001100111001111;
      // normal_words[17] = 32'b10010110110110111000001110100100;
      // normal_words[18] = 32'b01000011101000100010010010010101;
      // normal_words[19] = 32'b10110011110100100111110101111101;
      // normal_words[20] = 32'b11101011100010111101000111011001;
      // normal_words[21] = 32'b01100101001101001101111000001000;
      // normal_words[22] = 32'b01101110001101011010000000000100;
      // normal_words[23] = 32'b10011100010100110110111010101000;
      // normal_words[24] = 32'b11000100010001011110011001101111;
      // normal_words[25] = 32'b01101100011000011101111001010110;
      // normal_words[26] = 32'b11111011010001010001011000011011;
      // normal_words[27] = 32'b00111110111110101010100010010000;
      // normal_words[28] = 32'b11101011011010010011010101001001;
      // normal_words[29] = 32'b10001100100110010000001001111010;
      // normal_words[30] = 32'b01011000001111111111001101111100;
      // normal_words[31] = 32'b01100011011000111111100111010100;
      // normal_words[32] = 32'b11011100100010100011101001000100;
      // normal_words[33] = 32'b11111001100010011111110111110001;
      // normal_words[34] = 32'b01101011111000110001001011010110;
      // normal_words[35] = 32'b01011000110110101011111011000110;
      // normal_words[36] = 32'b00111011011100010001000100110010;
      // normal_words[37] = 32'b01100111110111001101001100001000;
      // normal_words[38] = 32'b11101010010101110000011000010101;
      // normal_words[39] = 32'b11111000000000110000110111000110;
      // normal_words[40] = 32'b11000111010110100000111111010110;
      // normal_words[41] = 32'b00001001101000001111000010101010;
      // normal_words[42] = 32'b01000111110100011010010001100010;
      // normal_words[43] = 32'b00100001101000111110101000000100;
      // normal_words[44] = 32'b00100101010111111000110000010101;
      // normal_words[45] = 32'b10111011010100110100010100011000;
      // normal_words[46] = 32'b10000100010111110101101111010100;
      // normal_words[47] = 32'b01011011110010001101110001011001;
      // normal_words[48] = 32'b10111010110111101000110001111001;
      // normal_words[49] = 32'b10101100000010111011011010100010;
      // normal_words[50] = 32'b01011100001110101000000101100100;
      // normal_words[51] = 32'b01010010100100011010111110111101;
      // normal_words[52] = 32'b01010111000001100010101110100100;
      // normal_words[53] = 32'b10000000110011101010101000001101;
      // normal_words[54] = 32'b01101011100100101011101110100110;
      // normal_words[55] = 32'b10101000101110001010110011100100;
      // normal_words[56] = 32'b11100100001111001011100101111110;
      // normal_words[57] = 32'b00010111110010111011101010100011;
      // normal_words[58] = 32'b00100011111111110110100110010001;
      // normal_words[59] = 32'b01101000110000111110101101011000;
      // normal_words[60] = 32'b10100100000001100100101011010111;
      // normal_words[61] = 32'b11001000101000110010100101111110;
      // normal_words[62] = 32'b01010110011110100110010011100001;
      // normal_words[63] = 32'b10111001000010001110110010100111;
      // normal_words[64] = 32'b10101001100101010111010001101111;
      // normal_words[65] = 32'b00110110001000010101011111100001;
      // normal_words[66] = 32'b10111101101000000100001110100010;
      // normal_words[67] = 32'b11011000101100001000000110111100;
      // normal_words[68] = 32'b10100011001001100111011110110101;
      // normal_words[69] = 32'b11111111111111010100100110110111;
      // normal_words[70] = 32'b10000101011011111111010000010111;
      // normal_words[71] = 32'b01100101110100101101100001111111;
      // normal_words[72] = 32'b11100011111011101010111110101011;
      // normal_words[73] = 32'b10011001101100110000011110011001;
      // normal_words[74] = 32'b11111001011011110011100010111100;
      // normal_words[75] = 32'b10010011011000101111111100000000;
      // normal_words[76] = 32'b10001111001010000001000010111011;
      // normal_words[77] = 32'b11101110100111000000100100010111;
      // normal_words[78] = 32'b00100110110100100101110011010111;
      // normal_words[79] = 32'b10110010110001111000000010111111;
      // normal_words[80] = 32'b11000100000000101001110010011100;
      // normal_words[81] = 32'b11111100011100100101001000111100;
      // normal_words[82] = 32'b11000010100100111110001111000001;
      // normal_words[83] = 32'b01100011111010000001111000111011;
      // normal_words[84] = 32'b11011110000011110001010111110111;
      // normal_words[85] = 32'b00110101011111011100011100100010;
      // normal_words[86] = 32'b11010011110100101001011001010100;
      // normal_words[87] = 32'b00101011110111011101010001101010;
      // normal_words[88] = 32'b10110111100111110111101101110000;
      // normal_words[89] = 32'b01000010001111000100010000100111;
      // normal_words[90] = 32'b00110100001001001010000101011011;
      // normal_words[91] = 32'b11001010100100101100010101001100;
      // normal_words[92] = 32'b11010011100011111000000100000011;
      // normal_words[93] = 32'b10101110000111100110010101011101;
      // normal_words[94] = 32'b00110001110000110100011110111101;
      // normal_words[95] = 32'b00011000111101000010010100001001;
      // normal_words[96] = 32'b00000110101001011101011110111110;
      // normal_words[97] = 32'b10000010100011001011000111110010;
      // normal_words[98] = 32'b10111111100001111001000111010010;
      // normal_words[99] = 32'b10000100000000001110001100100100;
      // normal_words[100] = 32'b10001101001110001101110000111111;
      // normal_words[101] = 32'b01101010011100001101001111111100;
      // normal_words[102] = 32'b01100010101101011100101010000000;
      // normal_words[103] = 32'b10111000010101111001111000101101;
      // normal_words[104] = 32'b11101010010110000100010111010111;
      // normal_words[105] = 32'b01010100111010111011011001100000;
      // normal_words[106] = 32'b00010110000110101100001010010101;
      // normal_words[107] = 32'b01111011101101110101101011111011;
      // normal_words[108] = 32'b00011001100110111000100000111110;
      // normal_words[109] = 32'b10110110001110010110100010001010;
      // normal_words[110] = 32'b00010101000110100010110001110111;
      // normal_words[111] = 32'b10001010001101110100010010100100;
      // normal_words[112] = 32'b00000001011111000011011010001001;
      // normal_words[113] = 32'b00011010011010111111011010011001;
      // normal_words[114] = 32'b10010001110101110011100001010100;
      // normal_words[115] = 32'b11111111110101100001001101011100;
      // normal_words[116] = 32'b11010101100011000110100001001101;
      // normal_words[117] = 32'b01000101010011000000101101010001;
      // normal_words[118] = 32'b01001101010101100000001010001111;
      // normal_words[119] = 32'b10101111110100011100010111110100;
      // normal_words[120] = 32'b01101000100100011101110001001101;
      // normal_words[121] = 32'b11000100011110111011001011011111;
      // normal_words[122] = 32'b01001011001001001100000001100011;
      // normal_words[123] = 32'b01010100011110001101100000101001;
      // normal_words[124] = 32'b11001100111010010101101111011010;
      // normal_words[125] = 32'b11111110011111110000110000100101;
      // normal_words[126] = 32'b11100000110111000001010111100100;
      // normal_words[127] = 32'b10001010000111100110011011000011;
      // normal_words[128] = 32'b11011110001111010111000010010111;
      // normal_words[129] = 32'b00011111001010001001001111100100;
      // normal_words[130] = 32'b10010011000101101000111000000100;
      // normal_words[131] = 32'b01010010110000101001110011011010;
      // normal_words[132] = 32'b00001101001110011000010100001111;
      // normal_words[133] = 32'b11000101111010010111110110001010;
      // normal_words[134] = 32'b00001011111110001111111100101000;
      // normal_words[135] = 32'b01000110000111000000101001101001;
      // normal_words[136] = 32'b01101100111010010110110011101011;
      // normal_words[137] = 32'b11101110110110011110101001010100;
      // normal_words[138] = 32'b11011100111001011000111001011111;
      // normal_words[139] = 32'b01001101000011110001101100010110;
      // normal_words[140] = 32'b10101000000100011100000100010101;
      // normal_words[141] = 32'b00010110011010010100100001010110;
      // normal_words[142] = 32'b00100100111111011000111101001001;
      // normal_words[143] = 32'b10000111001001100000000000001000;
      // normal_words[144] = 32'b10111000000111101001110010011101;
      // normal_words[145] = 32'b01110011101000011100010111001001;
      // normal_words[146] = 32'b10001110011000011101011000110010;
      // normal_words[147] = 32'b10101000001011110111010001001011;
      // normal_words[148] = 32'b11101011010111100010100000001101;
      // normal_words[149] = 32'b00001111001000011001101010100100;
      // normal_words[150] = 32'b11010000000000100011011101110111;
      // normal_words[151] = 32'b10000000110110011001110100110100;
      // normal_words[152] = 32'b00110111101001010101100100110110;
      // normal_words[153] = 32'b00111001001100000100010011110100;
      // normal_words[154] = 32'b01011101101011101110000111011101;
      // normal_words[155] = 32'b10001111011110011110011110111011;
      // normal_words[156] = 32'b11111001101101010110000101100000;
      // normal_words[157] = 32'b01101111000100011001010011011010;
      // normal_words[158] = 32'b10000011001001111100000111010111;
      // normal_words[159] = 32'b10001110011011010110101001110010;
      // normal_words[160] = 32'b01010001000111110110111010101000;
      // normal_words[161] = 32'b00000100110100001110101101100011;
      // normal_words[162] = 32'b10001111011010010010100000001111;
      // normal_words[163] = 32'b10101010011010100111001110111000;
      // normal_words[164] = 32'b01001110111011010001000000101001;
      // normal_words[165] = 32'b11011101000110101100000010101001;
      // normal_words[166] = 32'b11111001010010110011010001101001;
      // normal_words[167] = 32'b11001010011100110011011001110101;
      // normal_words[168] = 32'b10111110100001001100011110101001;
      // normal_words[169] = 32'b10000011011101111010010101100000;
      // normal_words[170] = 32'b10000110100101001001101111100111;
      // normal_words[171] = 32'b01001100000001100000011110010111;
      // normal_words[172] = 32'b11111101010101100010111101001000;
      // normal_words[173] = 32'b10000011111000110001110111110000;
      // normal_words[174] = 32'b10101101101111011100110001100101;
      // normal_words[175] = 32'b10011110010110010010100000001111;
      // normal_words[176] = 32'b00011011111011110011101001100010;
      // normal_words[177] = 32'b00100010001001011000010100111001;
      // normal_words[178] = 32'b00011001101111010010011101011001;
      // normal_words[179] = 32'b00000100011110001100100110011001;
      // normal_words[180] = 32'b11111000111101001110111111100100;
      // normal_words[181] = 32'b00111111001000011100101001100111;
      // normal_words[182] = 32'b10011011001001011001100001110111;
      // normal_words[183] = 32'b00010000100111000001010001101001;
      // normal_words[184] = 32'b01110110011001011110100110000111;
      // normal_words[185] = 32'b10111100101010100010101000000001;
      // normal_words[186] = 32'b11101100010101100101000011101110;
      // normal_words[187] = 32'b00100000110010100111011111110000;
      // normal_words[188] = 32'b10011110011010100010110110010011;
      // normal_words[189] = 32'b01101001000011110101100000110000;
      // normal_words[190] = 32'b11001111000001101100101010001100;
      // normal_words[191] = 32'b01010000010111111100111010011101;
      // normal_words[192] = 32'b00011010110110001100100000110100;
      // normal_words[193] = 32'b11111110110000000110100001110111;
      // normal_words[194] = 32'b11010011010001111011110101101110;
      // normal_words[195] = 32'b01010011010001110110100010110111;
      // normal_words[196] = 32'b01001101010011100101111101111000;
      // normal_words[197] = 32'b11111000100111110110110100001010;
      // normal_words[198] = 32'b10101111110101001000101011111110;
      // normal_words[199] = 32'b00000110011100010010100010110001;
      // normal_words[200] = 32'b00001100000001010110111001101001;
      // normal_words[201] = 32'b01100010001110110101011101000110;
      // normal_words[202] = 32'b01110101111111001011100011111110;
      // normal_words[203] = 32'b11001010011110101101100111010011;
      // normal_words[204] = 32'b00111100100011101011101000101110;
      // normal_words[205] = 32'b10011101100101100110101000111011;
      // normal_words[206] = 32'b11001010010001000111010110001000;
      // normal_words[207] = 32'b01001011001011010100111110000011;
      // normal_words[208] = 32'b00011110000010110111110010011010;
      // normal_words[209] = 32'b11000011101101110100001011011101;
      // normal_words[210] = 32'b10110010101100010100110110100111;
      // normal_words[211] = 32'b11110111011100001001010001111111;
      // normal_words[212] = 32'b01000100101000110011101110100111;
      // normal_words[213] = 32'b00001111100110000100101000111111;
      // normal_words[214] = 32'b11011011101011101000010001011010;
      // normal_words[215] = 32'b11111111000100001100101000011000;
      // normal_words[216] = 32'b01011111001010101100010100010010;
      // normal_words[217] = 32'b01110010111011001101010001001001;
      // normal_words[218] = 32'b11100000110111110111001110110000;
      // normal_words[219] = 32'b01000111011001110100111101001111;
      // normal_words[220] = 32'b11100011100101011001010110000000;
      // normal_words[221] = 32'b10000000001001101011101110111111;
      // normal_words[222] = 32'b01100101110011010101011100011100;
      // normal_words[223] = 32'b10001010000011110110001011011011;
      // normal_words[224] = 32'b11001010111000010000000001011110;
      // normal_words[225] = 32'b00011110000100000101010011100110;
      // normal_words[226] = 32'b11000000100010111101110100100001;
      // normal_words[227] = 32'b00101101101110010001110111110111;
      // normal_words[228] = 32'b01000001110000101101011100011100;
      // normal_words[229] = 32'b11101110010010001110011111000011;
      // normal_words[230] = 32'b11110010100101111110111001000010;
      // normal_words[231] = 32'b10000001001110100001000001001111;
      // normal_words[232] = 32'b10101101011100111100100100010010;
      // normal_words[233] = 32'b01001111100010011010001110010101;
      // normal_words[234] = 32'b00101100000101101000100111010110;
      // normal_words[235] = 32'b01000100011000000001101001001011;
      // normal_words[236] = 32'b01111011100001001001101100100101;
      // normal_words[237] = 32'b10011110101010101100111101010000;
      // normal_words[238] = 32'b10000000000000010011011001010010;
      // normal_words[239] = 32'b01100110000100001101110000101100;
      // normal_words[240] = 32'b10011110100100010001001100101100;
      // normal_words[241] = 32'b11001000101100011000010100011001;
      // normal_words[242] = 32'b00000011101000000111110110001101;
      // normal_words[243] = 32'b00111100100111101001001011110101;
      // normal_words[244] = 32'b01110110101100001010011101110001;
      // normal_words[245] = 32'b01000010100010011111010100001011;
      // normal_words[246] = 32'b00100001111100101100011000010001;
      // normal_words[247] = 32'b11110010001111010101011010010011;
      // normal_words[248] = 32'b01110010101100101110100011001110;
      // normal_words[249] = 32'b00110101011011001011100011011100;
      // normal_words[250] = 32'b10111100110000011110110101010111;
      // normal_words[251] = 32'b10000010011001111111111000000111;
      // normal_words[252] = 32'b00010011000111111111101100100000;
      // normal_words[253] = 32'b00111101110111101100110001100000;
      // normal_words[254] = 32'b00111101000100111011111110110011;
      // normal_words[255] = 32'b01011011011100100111101101001100;
      // normal_words[256] = 32'b11001001110010101101000101100111;
      // normal_words[257] = 32'b00011110001001011101010100100010;
      // normal_words[258] = 32'b00101010101111110000110011101010;
      // normal_words[259] = 32'b10000110101110011000110110111110;
      // normal_words[260] = 32'b01111100010001111110001101010000;
      // normal_words[261] = 32'b01111001101010000100101000000000;
      // normal_words[262] = 32'b00111010011101011011111001110110;
      // normal_words[263] = 32'b11111100110110111101000101000111;
      // normal_words[264] = 32'b00111010011100000100000111100111;
      // normal_words[265] = 32'b11001011110110111101100001000100;
      // normal_words[266] = 32'b11010100001010010011101100011010;
      // normal_words[267] = 32'b01101010010101100001011001001110;
      // normal_words[268] = 32'b01001001100010011010001001000000;
      // normal_words[269] = 32'b10101011011001111111110101001001;
      // normal_words[270] = 32'b01101001010000001100101101000111;
      // normal_words[271] = 32'b10111000000111000010110101100001;
      // normal_words[272] = 32'b01001110000011111000100101001110;
      // normal_words[273] = 32'b10111111000110110010001110111001;
      // normal_words[274] = 32'b11011010111010010010010111010011;
      // normal_words[275] = 32'b01110001101100010000100001000110;
      // normal_words[276] = 32'b10000100011011011101110100110111;
      // normal_words[277] = 32'b10011111011001001101001110011110;
      // normal_words[278] = 32'b01100011011111101010000110100010;
      // normal_words[279] = 32'b10010011011010001101101001000011;
      // normal_words[280] = 32'b11111100011010010101100001001001;
      // normal_words[281] = 32'b10011010001011101111011100111010;
      // normal_words[282] = 32'b11111000000101101000011010101101;
      // normal_words[283] = 32'b10110011111110010100010100110101;
      // normal_words[284] = 32'b10101000101111010011101101001010;
      // normal_words[285] = 32'b01100011100001010001110001110001;
      // normal_words[286] = 32'b11010011010111001001011010001100;
      // normal_words[287] = 32'b11000101110101100111101110011101;
      // normal_words[288] = 32'b00001011110001010011010111101001;
      // normal_words[289] = 32'b10011011101110110011110010100111;
      // normal_words[290] = 32'b01011100000110111111010000111001;
      // normal_words[291] = 32'b01110010110110101001100110110100;
      // normal_words[292] = 32'b01010101001111010001110100100011;
      // normal_words[293] = 32'b11111011101110001110001000101110;
      // normal_words[294] = 32'b01011010100000110111110010010011;
      // normal_words[295] = 32'b11111111100011101110011100010100;
      // normal_words[296] = 32'b11000101101010001000011011011111;
      // normal_words[297] = 32'b01010111001110111001001111011000;
      // normal_words[298] = 32'b11000001101110100101111001101000;
      // normal_words[299] = 32'b00011101101000101000000100001010;
      // normal_words[300] = 32'b10100001100011000000101110001100;
      // normal_words[301] = 32'b00101011000101110000000010101111;
      // normal_words[302] = 32'b11111111000000010001100101101001;
      // normal_words[303] = 32'b01000001001111001101111001010010;
      // normal_words[304] = 32'b01001010101110101100110011111101;
      // normal_words[305] = 32'b10011101001101000011011011101011;
      // normal_words[306] = 32'b00010100001011010011111101100100;
      // normal_words[307] = 32'b10111100111011001000011010100111;
      // normal_words[308] = 32'b00100000000001000010111010010100;
      // normal_words[309] = 32'b01100110110110000100011110110011;
      // normal_words[310] = 32'b10110110110011101001001010101110;
      // normal_words[311] = 32'b10000110110100101111111011010010;
      // normal_words[312] = 32'b11001110001110110100011010101001;
      // normal_words[313] = 32'b01000111101000101110010010001000;
      // normal_words[314] = 32'b01110011110011101101111110011101;
      // normal_words[315] = 32'b10101100010111011000000111110001;
      // normal_words[316] = 32'b10001111100100101010000111010010;
      // normal_words[317] = 32'b10111110111101011011101100110010;
      // normal_words[318] = 32'b00110101110100000111011001110100;
      // normal_words[319] = 32'b10110001110111010010011000100110;
      // normal_words[320] = 32'b11101111100000110100100010000110;
      // normal_words[321] = 32'b10011001000101111001100010010110;
      // normal_words[322] = 32'b00111010001101111111010000110001;
      // normal_words[323] = 32'b10000011001100010101011001100101;
      // normal_words[324] = 32'b10110000111010101100000001101110;
      // normal_words[325] = 32'b01101000001111100111011101110011;
      // normal_words[326] = 32'b01000000101111011010110111100010;
      // normal_words[327] = 32'b10100010100100111100110000111110;
      // normal_words[328] = 32'b11101111000101001001011111100001;
      // normal_words[329] = 32'b00100101100011000110001100111001;
      // normal_words[330] = 32'b11101000000001010011111110101111;
      // normal_words[331] = 32'b11000011110001100100100010001001;
      // normal_words[332] = 32'b10110100101101001111000010100011;
      // normal_words[333] = 32'b01100101111110101110000100001101;
      // normal_words[334] = 32'b01011011000001001110001010100111;
      // normal_words[335] = 32'b01000001101111001010010110110010;
      // normal_words[336] = 32'b10001010010011010000101010111000;
      // normal_words[337] = 32'b11101000011011010111000010011111;
      // normal_words[338] = 32'b00011100011101101110111100100101;
      // normal_words[339] = 32'b11000000000101000011101110111010;
      // normal_words[340] = 32'b10001111000001001001111110011011;
      // normal_words[341] = 32'b00110101110111011110110001000010;
      // normal_words[342] = 32'b10111111000101001100100111001111;
      // normal_words[343] = 32'b10001110110101101111011100100111;
      // normal_words[344] = 32'b00001100111000010000001000011101;
      // normal_words[345] = 32'b10001000011000001111010111001111;
      // normal_words[346] = 32'b11000001110110100111101100001010;
      // normal_words[347] = 32'b01100101110001111001100110011001;
      // normal_words[348] = 32'b00110011111101101000000000011101;
      // normal_words[349] = 32'b10110100101100111111010101110011;
      // normal_words[350] = 32'b10001101001011000011111111100111;
      // normal_words[351] = 32'b00010000101100011111111010011000;
      // normal_words[352] = 32'b11110111010111010100111100011001;
      // normal_words[353] = 32'b10110010111000100010001100111000;
      // normal_words[354] = 32'b00101100110100101101010111111100;
      // normal_words[355] = 32'b00100111100011011011101011011001;
      // normal_words[356] = 32'b00110000011100110000011000010101;
      // normal_words[357] = 32'b11111001111000010011000011000011;
      // normal_words[358] = 32'b10101010010100000010111000100110;
      // normal_words[359] = 32'b00110111111100111001001010110011;
      // normal_words[360] = 32'b11000001101010000001001100000101;
      // normal_words[361] = 32'b01110100100111111001011101101001;
      // normal_words[362] = 32'b11101110100000001011001110111001;
      // normal_words[363] = 32'b00101000110101001110111001001100;
      // normal_words[364] = 32'b00101001111100000101101111110101;
      // normal_words[365] = 32'b00000010101001100001010100000010;
      // normal_words[366] = 32'b01110000001100010110110101010100;
      // normal_words[367] = 32'b01011010101110101001100101110110;
      // normal_words[368] = 32'b11001101010001100100001110011011;
      // normal_words[369] = 32'b01110101100100101010110110011110;
      // normal_words[370] = 32'b00000011100101010011001111000001;
      // normal_words[371] = 32'b00111110010101111011000110100010;
      // normal_words[372] = 32'b01001100100001000011101110000100;
      // normal_words[373] = 32'b00110000100100010101000110110100;
      // normal_words[374] = 32'b11100111110110111100011100000010;
      // normal_words[375] = 32'b01110101110000111011000000101101;
      // normal_words[376] = 32'b11101110001010011101001111000111;
      // normal_words[377] = 32'b11011111100011001110010110100110;
      // normal_words[378] = 32'b10011001001111001100100000111101;
      // normal_words[379] = 32'b00011101011011011111101001001111;
      // normal_words[380] = 32'b01001010101010000001110111000100;
      // normal_words[381] = 32'b01110000010100100000010010101000;
      // normal_words[382] = 32'b10100101000011101001110000010100;
      // normal_words[383] = 32'b11010110010111101011011001010110;
      // normal_words[384] = 32'b11100011110011100001110010101110;
      // normal_words[385] = 32'b01101101001011010011011100111101;
      // normal_words[386] = 32'b11101100010001011101010101010101;
      // normal_words[387] = 32'b11101110000100001001000000001100;
      // normal_words[388] = 32'b01111101100100100001111100011001;
      // normal_words[389] = 32'b11000001011111000101011000101011;
      // normal_words[390] = 32'b00011101100011111010010100001001;
      // normal_words[391] = 32'b01101011010010101110011000000001;
      // normal_words[392] = 32'b01000100011011111101111111000100;
      // normal_words[393] = 32'b11100111100110001110101100111111;
      // normal_words[394] = 32'b01001001100101101101001101001101;
      // normal_words[395] = 32'b11100000001101110111101001111000;
      // normal_words[396] = 32'b01110111001010001001010101101110;
      // normal_words[397] = 32'b11111010011100001110000100100101;
      // normal_words[398] = 32'b01101011110010100100100110011000;
      // normal_words[399] = 32'b10011101110101100010011000101110;
      // normal_words[400] = 32'b00011110101000100101011011011101;
      // normal_words[401] = 32'b11000001111000000000110110101110;
      // normal_words[402] = 32'b00111110100110001100010011110100;
      // normal_words[403] = 32'b01010101011101110100100000110010;
      // normal_words[404] = 32'b10110001101001110011001110011101;
      // normal_words[405] = 32'b11000111101010010111101010101001;
      // normal_words[406] = 32'b01111100000001001011010010001010;
      // normal_words[407] = 32'b00011011001000100000011110011111;
      // normal_words[408] = 32'b10001100010101101011100001010110;
      // normal_words[409] = 32'b11100111111010010010000111101110;
      // normal_words[410] = 32'b01101110011100111111111001001110;
      // normal_words[411] = 32'b11101010011111111110010101010110;
      // normal_words[412] = 32'b01001000100010100010010111000000;
      // normal_words[413] = 32'b00000011001010111111100111100000;
      // normal_words[414] = 32'b01111010011101101001111000110110;
      // normal_words[415] = 32'b00000100011000010011101110101000;
      // normal_words[416] = 32'b00100100000100000111011100001011;
      // normal_words[417] = 32'b00001001011100011110011100000011;
      // normal_words[418] = 32'b10101100011110010000011010011001;
      // normal_words[419] = 32'b01101100100001001000111000001011;
      // normal_words[420] = 32'b00101011010000100110000001110101;
      // normal_words[421] = 32'b00001001111000100110011110110001;
      // normal_words[422] = 32'b10111100110011100110100110110111;
      // normal_words[423] = 32'b11010111110000010011101010110011;
      // normal_words[424] = 32'b10100011111010000111100000010001;
      // normal_words[425] = 32'b01010110010011110100001101011011;
      // normal_words[426] = 32'b01011000001000101111101101100100;
      // normal_words[427] = 32'b10110001100110010000100001001110;
      // normal_words[428] = 32'b00111010110001100100001001100000;
      // normal_words[429] = 32'b11111010001110100111100100000101;
      // normal_words[430] = 32'b10001001011000111101100010000101;
      // normal_words[431] = 32'b11101101101110111011001001100001;
      // normal_words[432] = 32'b11100011000111000011011111001011;
      // normal_words[433] = 32'b10010001101111100010111010010001;
      // normal_words[434] = 32'b00101100011010011110110100110111;
      // normal_words[435] = 32'b11111110001010111011100110011010;
      // normal_words[436] = 32'b00110101011110100010100110100101;
      // normal_words[437] = 32'b01000101011111100100100110011111;
      // normal_words[438] = 32'b01010100001101111001110111111001;
      // normal_words[439] = 32'b10101010011101110000110010011011;
      // normal_words[440] = 32'b01110001011000000111000110110100;
      // normal_words[441] = 32'b10101110101000110111010100001111;
      // normal_words[442] = 32'b01000111110001001111000010100100;
      // normal_words[443] = 32'b10000101011111101110111110111101;
      // normal_words[444] = 32'b01111000001001111110010011111011;
      // normal_words[445] = 32'b11001001010110011010101110001100;
      // normal_words[446] = 32'b10100110000001010011011101011101;
      // normal_words[447] = 32'b10010000010100010010100000000011;
      // normal_words[448] = 32'b11100111000001001110011001011011;
      // normal_words[449] = 32'b00111010000100001001000100111110;
      // normal_words[450] = 32'b10110010100101011100101101010001;
      // normal_words[451] = 32'b10110011011000001101001101110110;
      // normal_words[452] = 32'b01010000000001000100100111000011;
      // normal_words[453] = 32'b11001100010110010111011110110111;
      // normal_words[454] = 32'b10100000011110011001111110010110;
      // normal_words[455] = 32'b11001111100110111101001000001011;
      // normal_words[456] = 32'b01000100111100110111110100101101;
      // normal_words[457] = 32'b00100010101110001100110100010010;
      // normal_words[458] = 32'b10110100110000000000101101010000;
      // normal_words[459] = 32'b00011001100100100000110001010111;
      // normal_words[460] = 32'b00000011000110001001010011100000;
      // normal_words[461] = 32'b00000111001011001010110110011101;
      // normal_words[462] = 32'b01010000110000100011000010000001;
      // normal_words[463] = 32'b11011011001000011010110110010000;
      // normal_words[464] = 32'b10000110001101010111011101011011;
      // normal_words[465] = 32'b11111111000011110101010100100000;
      // normal_words[466] = 32'b01000010011111100010101110001001;
      // normal_words[467] = 32'b00110011010111011101010000101110;
      // normal_words[468] = 32'b00000111101011010111011000010111;
      // normal_words[469] = 32'b00000110101101010100100100111100;
      // normal_words[470] = 32'b01111110101010010110000110111000;
      // normal_words[471] = 32'b10111101010011101011100000101011;
      // normal_words[472] = 32'b00110001010111110111100101001110;
      // normal_words[473] = 32'b10111110010001011000000011000011;
      // normal_words[474] = 32'b00011101001011011000011011100110;
      // normal_words[475] = 32'b10011111111010001001101101111011;
      // normal_words[476] = 32'b10101111110011011000010100001111;
      // normal_words[477] = 32'b11100000000100110111110000101000;
      // normal_words[478] = 32'b11000000111111010000000001001001;
      // normal_words[479] = 32'b01010000011000101101010000000000;
      // normal_words[480] = 32'b00110011100010111001100010101100;
      // normal_words[481] = 32'b10011101000111111001001000010010;
      // normal_words[482] = 32'b01101000110110101010110111110001;
      // normal_words[483] = 32'b00010011010111110110111111000111;
      // normal_words[484] = 32'b10000001001011001100101010100000;
      // normal_words[485] = 32'b11010111010000000000110111111010;
      // normal_words[486] = 32'b00100011111110010010111110000101;
      // normal_words[487] = 32'b10110110110100111101111001000111;
      // normal_words[488] = 32'b01000110101010111110110111000010;
      // normal_words[489] = 32'b10000001001011101110010101110011;
      // normal_words[490] = 32'b10100001100011001100100000110101;
      // normal_words[491] = 32'b01000110110001011001110110010111;
      // normal_words[492] = 32'b00101010100101000100010110010011;
      // normal_words[493] = 32'b01101010000010110111011100110110;
      // normal_words[494] = 32'b10010110000100111001010110100011;
      // normal_words[495] = 32'b01011110110110000101000010001110;
      // normal_words[496] = 32'b11011110101010100110001111110110;
      // normal_words[497] = 32'b01111100100110111110111011000101;
      // normal_words[498] = 32'b11101111001100111101011100001101;
      // normal_words[499] = 32'b10010110000000100110010110101111;
      // normal_words[500] = 32'b01101010110010001010100001110100;
      // normal_words[501] = 32'b00011110000101110101100111101111;
      // normal_words[502] = 32'b11101111001011110010101110100000;
      // normal_words[503] = 32'b10000010000111101001000100111000;
      // normal_words[504] = 32'b00000011111000000010011110011110;
      // normal_words[505] = 32'b10011110010000111101001010000100;
      // normal_words[506] = 32'b00110101101011010100110100011010;
      // normal_words[507] = 32'b00110010100011100111100101100010;
      // normal_words[508] = 32'b01111101011010000001100011110101;
      // normal_words[509] = 32'b11001100111100001001000101011000;
      // normal_words[510] = 32'b00111100011010110001110110110011;
      // normal_words[511] = 32'b01100101100000101100110101001101;
      // normal_words[512] = 32'b10011100100010000001100000100001;
      // normal_words[513] = 32'b00000100101000100000000011101011;
      // normal_words[514] = 32'b10010100100110101110111101011101;
      // normal_words[515] = 32'b01011001011111000011111111011010;
      // normal_words[516] = 32'b11010100100100101011011010101001;
      // normal_words[517] = 32'b01100101000110010000011000010010;
      // normal_words[518] = 32'b01011011101111110100111110101110;
      // normal_words[519] = 32'b10000000011010100011001111011000;
      // normal_words[520] = 32'b11011111111001000001101010000111;
      // normal_words[521] = 32'b00011101100000010010000000001010;
      // normal_words[522] = 32'b00110011111100011111110101001111;
      // normal_words[523] = 32'b10010000111001010110110000011101;
      // normal_words[524] = 32'b10101011000100101100011011000010;
      // normal_words[525] = 32'b10111000110110010101110011110001;
      // normal_words[526] = 32'b01101011100111000011010010000101;
      // normal_words[527] = 32'b10110100101001111100100000010001;
      // normal_words[528] = 32'b00101111100111111101111010111011;
      // normal_words[529] = 32'b00111100000101000011011000100101;
      // normal_words[530] = 32'b11101010111111100110001000010101;
      // normal_words[531] = 32'b11001101011010011010111000110000;
      // normal_words[532] = 32'b10101110000100111110111000110010;
      // normal_words[533] = 32'b11011100011101111001001110000010;
      // normal_words[534] = 32'b00011101100001101001001001111101;
      // normal_words[535] = 32'b01000001110101101101000111101111;
      // normal_words[536] = 32'b11101010000111101001101010011001;
      // normal_words[537] = 32'b11010100000101010000000011110111;
      // normal_words[538] = 32'b01001110101111011010011101000111;
      // normal_words[539] = 32'b01001001001000010001001101101001;
      // normal_words[540] = 32'b10110100001100010000111111000101;
      // normal_words[541] = 32'b11000001100011111110001110110001;
      // normal_words[542] = 32'b01001111100000101000110001110110;
      // normal_words[543] = 32'b00101011100001100100111001101110;
      // normal_words[544] = 32'b11011001111000001101111100101101;
      // normal_words[545] = 32'b01111000101100011010000101001101;
      // normal_words[546] = 32'b10111001000011100011011111111110;
      // normal_words[547] = 32'b00001111001111110101001111100111;
      // normal_words[548] = 32'b01100010001001111000100111111101;
      // normal_words[549] = 32'b01010101001100001011010001101110;
      // normal_words[550] = 32'b01100100010110100000011110011111;
      // normal_words[551] = 32'b01010111011111010111100010001011;
      // normal_words[552] = 32'b00000000000000000000000000000101;


      // for (j = 0; j < WEIGHT; j = j + 1) begin
      //    encrypt_index(sparse_pairs[j], j);  // sparse_pairs[i]를 TEXTIN으로 사용, key 값은 i (0~65)
      // end

      // for (j =WEIGHT; j < MEM_SIZE + WEIGHT; j = j + 1) begin
      //    encrypt_text(normal_words[j - WEIGHT], j);  // normal_words[i-66]를 TEXTIN으로 사용, key 값은 i (66~618)
      // end

      // $display("done!");
      // #(pUSB_CLOCK_PERIOD*10);
      // if (errors)
      //    $display("SIMULATION FAILED (%0d errors, %0d warnings).", errors, warnings);
      // else
      //    $display("Simulation passed (%0d warnings).", warnings);
      // $finish;

   end

   // maintain a cycle counter
   always @(posedge clk) begin
      if (pushbutton == 0)
         cycle <= 0;
      else
         cycle <= cycle + 1;
   end


   // timeout thread:
   initial begin
      #(pUSB_CLOCK_PERIOD*pTIMEOUT);
      errors = errors + 1;
      $display("ERROR: global timeout");
      $display("SIMULATION FAILED (%0d errors).", errors);
      $finish;
   end


   reg read_select;

   assign usb_data = read_select? 8'bz : usb_wdata;
   assign tio_clkin = pll_clk1;

   always @(*) begin
      if (usb_wrn == 1'b0)
         read_select = 1'b0;
      else if (usb_rdn == 1'b0)
         read_select = 1'b1;
   end


   always #(pUSB_CLOCK_PERIOD/2) usb_clk = !usb_clk;
   always #(pPLL_CLOCK_PERIOD/2) pll_clk1 = !pll_clk1;

   wire #1 usb_rdn_out = usb_rdn;
   wire #1 usb_wrn_out = usb_wrn;
   wire #1 usb_cen_out = usb_cen;
   wire #1 usb_trigger_out = usb_trigger;

   wire trigger; // TODO: use it?

   cw305_top #(
      .pBYTECNT_SIZE            (pBYTECNT_SIZE),
      .pADDR_WIDTH              (pADDR_WIDTH)
   ) U_dut (
      .usb_clk                  (usb_clk & usb_clk_enable),
      .usb_data                 (usb_data),
      .usb_addr                 (usb_addr),
      .usb_rdn                  (usb_rdn_out),
      .usb_wrn                  (usb_wrn_out),
      .usb_cen                  (usb_cen_out),
      .usb_trigger              (usb_trigger_out),
      .j16_sel                  (j16_sel),
      .k16_sel                  (k16_sel),
      .k15_sel                  (k15_sel),
      .l14_sel                  (l14_sel),
      .pushbutton               (pushbutton),
      .led1                     (led1),
      .led2                     (led2),
      .led3                     (led3),
      .pll_clk1                 (pll_clk1),
      .tio_trigger              (trigger),
      .tio_clkout               (),             // unused
      .tio_clkin                (tio_clkin)
   );


   task wait_done;
      reg busy;
      begin
         busy = 1;
         while (busy == 1) begin
            //$display("checking busy...");
            read_byte(0, `REG_CRYPT_GO, 0, busy);
         end
      end
   endtask


endmodule

`default_nettype wire

